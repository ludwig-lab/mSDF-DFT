-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 12 2024 10:20:51

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "top_test" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of top_test
entity top_test is
port (
    o_X : out std_logic_vector(31 downto 0);
    i_ref_clk : in std_logic;
    done : out std_logic;
    i_rst : in std_logic);
end top_test;

-- Architecture of top_test
-- View name is \INTERFACE\
architecture \INTERFACE\ of top_test is

signal \N__7068\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7041\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7023\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7014\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7005\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7003\ : std_logic;
signal \N__6996\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6994\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6986\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6978\ : std_logic;
signal \N__6977\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6969\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6959\ : std_logic;
signal \N__6958\ : std_logic;
signal \N__6951\ : std_logic;
signal \N__6950\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6941\ : std_logic;
signal \N__6940\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6923\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6915\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6906\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6904\ : std_logic;
signal \N__6897\ : std_logic;
signal \N__6896\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6888\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6879\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6877\ : std_logic;
signal \N__6870\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6868\ : std_logic;
signal \N__6861\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6859\ : std_logic;
signal \N__6852\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6850\ : std_logic;
signal \N__6843\ : std_logic;
signal \N__6842\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6832\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6824\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6816\ : std_logic;
signal \N__6815\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6807\ : std_logic;
signal \N__6806\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6797\ : std_logic;
signal \N__6796\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6788\ : std_logic;
signal \N__6787\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6771\ : std_logic;
signal \N__6770\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6731\ : std_logic;
signal \N__6728\ : std_logic;
signal \N__6725\ : std_logic;
signal \N__6722\ : std_logic;
signal \N__6719\ : std_logic;
signal \N__6716\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6710\ : std_logic;
signal \N__6707\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6701\ : std_logic;
signal \N__6698\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6696\ : std_logic;
signal \N__6695\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6689\ : std_logic;
signal \N__6686\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6649\ : std_logic;
signal \N__6646\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6632\ : std_logic;
signal \N__6629\ : std_logic;
signal \N__6626\ : std_logic;
signal \N__6623\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6608\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6602\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6596\ : std_logic;
signal \N__6593\ : std_logic;
signal \N__6590\ : std_logic;
signal \N__6587\ : std_logic;
signal \N__6584\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6579\ : std_logic;
signal \N__6578\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6576\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6574\ : std_logic;
signal \N__6573\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6571\ : std_logic;
signal \N__6570\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6568\ : std_logic;
signal \N__6567\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6533\ : std_logic;
signal \N__6530\ : std_logic;
signal \N__6529\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6519\ : std_logic;
signal \N__6518\ : std_logic;
signal \N__6517\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6515\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6513\ : std_logic;
signal \N__6512\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6510\ : std_logic;
signal \N__6509\ : std_logic;
signal \N__6508\ : std_logic;
signal \N__6507\ : std_logic;
signal \N__6506\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6503\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6495\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6491\ : std_logic;
signal \N__6490\ : std_logic;
signal \N__6487\ : std_logic;
signal \N__6484\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6371\ : std_logic;
signal \N__6368\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6344\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6332\ : std_logic;
signal \N__6329\ : std_logic;
signal \N__6326\ : std_logic;
signal \N__6323\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6314\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6308\ : std_logic;
signal \N__6305\ : std_logic;
signal \N__6302\ : std_logic;
signal \N__6299\ : std_logic;
signal \N__6296\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6287\ : std_logic;
signal \N__6284\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6278\ : std_logic;
signal \N__6275\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6263\ : std_logic;
signal \N__6260\ : std_logic;
signal \N__6257\ : std_logic;
signal \N__6254\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6242\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6233\ : std_logic;
signal \N__6230\ : std_logic;
signal \N__6227\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6203\ : std_logic;
signal \N__6200\ : std_logic;
signal \N__6197\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6182\ : std_logic;
signal \N__6179\ : std_logic;
signal \N__6176\ : std_logic;
signal \N__6173\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6155\ : std_logic;
signal \N__6152\ : std_logic;
signal \N__6149\ : std_logic;
signal \N__6146\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6139\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6133\ : std_logic;
signal \N__6130\ : std_logic;
signal \N__6127\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6121\ : std_logic;
signal \N__6116\ : std_logic;
signal \N__6113\ : std_logic;
signal \N__6110\ : std_logic;
signal \N__6107\ : std_logic;
signal \N__6104\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6098\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6077\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6062\ : std_logic;
signal \N__6059\ : std_logic;
signal \N__6056\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6041\ : std_logic;
signal \N__6038\ : std_logic;
signal \N__6035\ : std_logic;
signal \N__6034\ : std_logic;
signal \N__6033\ : std_logic;
signal \N__6032\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6027\ : std_logic;
signal \N__6026\ : std_logic;
signal \N__6023\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6002\ : std_logic;
signal \N__5997\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5984\ : std_logic;
signal \N__5969\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5963\ : std_logic;
signal \N__5960\ : std_logic;
signal \N__5957\ : std_logic;
signal \N__5954\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5952\ : std_logic;
signal \N__5951\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5945\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5942\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5936\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5934\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5931\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5928\ : std_logic;
signal \N__5927\ : std_logic;
signal \N__5926\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5922\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5901\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5898\ : std_logic;
signal \N__5897\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5894\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5891\ : std_logic;
signal \N__5890\ : std_logic;
signal \N__5889\ : std_logic;
signal \N__5888\ : std_logic;
signal \N__5887\ : std_logic;
signal \N__5886\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5881\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5873\ : std_logic;
signal \N__5872\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5869\ : std_logic;
signal \N__5868\ : std_logic;
signal \N__5865\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5840\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5836\ : std_logic;
signal \N__5835\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5826\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5791\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5759\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5740\ : std_logic;
signal \N__5723\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5699\ : std_logic;
signal \N__5696\ : std_logic;
signal \N__5693\ : std_logic;
signal \N__5690\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5686\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5663\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5622\ : std_logic;
signal \N__5619\ : std_logic;
signal \N__5616\ : std_logic;
signal \N__5609\ : std_logic;
signal \N__5606\ : std_logic;
signal \N__5601\ : std_logic;
signal \N__5596\ : std_logic;
signal \N__5593\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5582\ : std_logic;
signal \N__5579\ : std_logic;
signal \N__5576\ : std_logic;
signal \N__5573\ : std_logic;
signal \N__5570\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5552\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5543\ : std_logic;
signal \N__5540\ : std_logic;
signal \N__5537\ : std_logic;
signal \N__5534\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5528\ : std_logic;
signal \N__5525\ : std_logic;
signal \N__5522\ : std_logic;
signal \N__5519\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5492\ : std_logic;
signal \N__5489\ : std_logic;
signal \N__5486\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5480\ : std_logic;
signal \N__5477\ : std_logic;
signal \N__5474\ : std_logic;
signal \N__5471\ : std_logic;
signal \N__5468\ : std_logic;
signal \N__5465\ : std_logic;
signal \N__5462\ : std_logic;
signal \N__5459\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5453\ : std_logic;
signal \N__5450\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5441\ : std_logic;
signal \N__5438\ : std_logic;
signal \N__5435\ : std_logic;
signal \N__5432\ : std_logic;
signal \N__5429\ : std_logic;
signal \N__5426\ : std_logic;
signal \N__5423\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5411\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5396\ : std_logic;
signal \N__5393\ : std_logic;
signal \N__5390\ : std_logic;
signal \N__5387\ : std_logic;
signal \N__5384\ : std_logic;
signal \N__5381\ : std_logic;
signal \N__5378\ : std_logic;
signal \N__5375\ : std_logic;
signal \N__5372\ : std_logic;
signal \N__5369\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5360\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5348\ : std_logic;
signal \N__5345\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5338\ : std_logic;
signal \N__5335\ : std_logic;
signal \N__5332\ : std_logic;
signal \N__5329\ : std_logic;
signal \N__5324\ : std_logic;
signal \N__5323\ : std_logic;
signal \N__5320\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5308\ : std_logic;
signal \N__5305\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5288\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5279\ : std_logic;
signal \N__5276\ : std_logic;
signal \N__5273\ : std_logic;
signal \N__5270\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5252\ : std_logic;
signal \N__5249\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5211\ : std_logic;
signal \N__5208\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5201\ : std_logic;
signal \N__5198\ : std_logic;
signal \N__5195\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5180\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5167\ : std_logic;
signal \N__5166\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5141\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5122\ : std_logic;
signal \N__5119\ : std_logic;
signal \N__5116\ : std_logic;
signal \N__5111\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5091\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5076\ : std_logic;
signal \N__5073\ : std_logic;
signal \N__5072\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5066\ : std_logic;
signal \N__5065\ : std_logic;
signal \N__5062\ : std_logic;
signal \N__5059\ : std_logic;
signal \N__5056\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5027\ : std_logic;
signal \N__5024\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5018\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5000\ : std_logic;
signal \N__4997\ : std_logic;
signal \N__4994\ : std_logic;
signal \N__4991\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4985\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4976\ : std_logic;
signal \N__4975\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4960\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4955\ : std_logic;
signal \N__4952\ : std_logic;
signal \N__4949\ : std_logic;
signal \N__4946\ : std_logic;
signal \N__4939\ : std_logic;
signal \N__4938\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4905\ : std_logic;
signal \N__4902\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4892\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4886\ : std_logic;
signal \N__4883\ : std_logic;
signal \N__4880\ : std_logic;
signal \N__4877\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4835\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4814\ : std_logic;
signal \N__4811\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4772\ : std_logic;
signal \N__4769\ : std_logic;
signal \N__4766\ : std_logic;
signal \N__4763\ : std_logic;
signal \N__4762\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4755\ : std_logic;
signal \N__4752\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4750\ : std_logic;
signal \N__4747\ : std_logic;
signal \N__4744\ : std_logic;
signal \N__4741\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4735\ : std_logic;
signal \N__4732\ : std_logic;
signal \N__4725\ : std_logic;
signal \N__4722\ : std_logic;
signal \N__4719\ : std_logic;
signal \N__4716\ : std_logic;
signal \N__4713\ : std_logic;
signal \N__4706\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4699\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4682\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4675\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4664\ : std_logic;
signal \N__4661\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4657\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4646\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4634\ : std_logic;
signal \N__4633\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4622\ : std_logic;
signal \N__4619\ : std_logic;
signal \N__4616\ : std_logic;
signal \N__4613\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4601\ : std_logic;
signal \N__4598\ : std_logic;
signal \N__4595\ : std_logic;
signal \N__4592\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4586\ : std_logic;
signal \N__4583\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4565\ : std_logic;
signal \N__4562\ : std_logic;
signal \N__4559\ : std_logic;
signal \N__4556\ : std_logic;
signal \N__4553\ : std_logic;
signal \N__4550\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4538\ : std_logic;
signal \N__4535\ : std_logic;
signal \N__4532\ : std_logic;
signal \N__4529\ : std_logic;
signal \N__4526\ : std_logic;
signal \N__4523\ : std_logic;
signal \N__4520\ : std_logic;
signal \N__4517\ : std_logic;
signal \N__4514\ : std_logic;
signal \N__4511\ : std_logic;
signal \N__4508\ : std_logic;
signal \N__4505\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4484\ : std_logic;
signal \N__4481\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4445\ : std_logic;
signal \N__4442\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4436\ : std_logic;
signal \N__4433\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4403\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4394\ : std_logic;
signal \N__4391\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4379\ : std_logic;
signal \N__4376\ : std_logic;
signal \N__4373\ : std_logic;
signal \N__4370\ : std_logic;
signal \N__4367\ : std_logic;
signal \N__4364\ : std_logic;
signal \N__4361\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4349\ : std_logic;
signal \N__4346\ : std_logic;
signal \N__4343\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4307\ : std_logic;
signal \N__4304\ : std_logic;
signal \N__4301\ : std_logic;
signal \N__4298\ : std_logic;
signal \N__4295\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4265\ : std_logic;
signal \N__4262\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4247\ : std_logic;
signal \N__4244\ : std_logic;
signal \N__4241\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4235\ : std_logic;
signal \N__4232\ : std_logic;
signal \N__4229\ : std_logic;
signal \N__4226\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4222\ : std_logic;
signal \N__4219\ : std_logic;
signal \N__4216\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4208\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4202\ : std_logic;
signal \N__4199\ : std_logic;
signal \N__4196\ : std_logic;
signal \N__4193\ : std_logic;
signal \N__4190\ : std_logic;
signal \N__4187\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4181\ : std_logic;
signal \N__4178\ : std_logic;
signal \N__4175\ : std_logic;
signal \N__4172\ : std_logic;
signal \N__4169\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4163\ : std_logic;
signal \N__4160\ : std_logic;
signal \N__4157\ : std_logic;
signal \N__4154\ : std_logic;
signal \N__4151\ : std_logic;
signal \N__4148\ : std_logic;
signal \N__4145\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4133\ : std_logic;
signal \N__4130\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4115\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4007\ : std_logic;
signal \N__4004\ : std_logic;
signal \N__4001\ : std_logic;
signal \N__3998\ : std_logic;
signal \N__3995\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3983\ : std_logic;
signal \N__3980\ : std_logic;
signal \N__3977\ : std_logic;
signal \N__3974\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3962\ : std_logic;
signal \N__3959\ : std_logic;
signal \N__3956\ : std_logic;
signal \N__3953\ : std_logic;
signal \N__3950\ : std_logic;
signal \N__3947\ : std_logic;
signal \N__3944\ : std_logic;
signal \N__3941\ : std_logic;
signal \N__3938\ : std_logic;
signal \N__3935\ : std_logic;
signal \N__3932\ : std_logic;
signal \N__3929\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3917\ : std_logic;
signal \N__3914\ : std_logic;
signal \N__3911\ : std_logic;
signal \N__3908\ : std_logic;
signal \N__3905\ : std_logic;
signal \N__3902\ : std_logic;
signal \N__3899\ : std_logic;
signal \N__3896\ : std_logic;
signal \N__3893\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3887\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3881\ : std_logic;
signal \N__3878\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3854\ : std_logic;
signal \N__3851\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3818\ : std_logic;
signal \N__3815\ : std_logic;
signal \N__3812\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3767\ : std_logic;
signal \N__3764\ : std_logic;
signal \N__3761\ : std_logic;
signal \N__3758\ : std_logic;
signal \N__3755\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3713\ : std_logic;
signal \N__3710\ : std_logic;
signal \N__3707\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3698\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3683\ : std_logic;
signal \N__3680\ : std_logic;
signal \N__3677\ : std_logic;
signal \N__3674\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3668\ : std_logic;
signal \N__3665\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3647\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3641\ : std_logic;
signal \N__3638\ : std_logic;
signal \N__3635\ : std_logic;
signal \N__3632\ : std_logic;
signal \N__3629\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3620\ : std_logic;
signal \N__3617\ : std_logic;
signal \N__3614\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3596\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3539\ : std_logic;
signal \N__3536\ : std_logic;
signal \N__3533\ : std_logic;
signal \N__3530\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3521\ : std_logic;
signal \N__3518\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3505\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3501\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3485\ : std_logic;
signal \N__3482\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3431\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3422\ : std_logic;
signal \N__3419\ : std_logic;
signal \N__3416\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3407\ : std_logic;
signal \N__3404\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3392\ : std_logic;
signal \N__3389\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3368\ : std_logic;
signal \N__3365\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3362\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3360\ : std_logic;
signal \N__3359\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3357\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3354\ : std_logic;
signal \N__3353\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3350\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3347\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3344\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3342\ : std_logic;
signal \N__3341\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3339\ : std_logic;
signal \N__3338\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3278\ : std_logic;
signal \N__3275\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3266\ : std_logic;
signal sys_clk_g : std_logic;
signal sys_clk : std_logic;
signal \GNDG0\ : std_logic;
signal i_ref_clk_c : std_logic;
signal \VCCG0\ : std_logic;
signal i_rst_c_i : std_logic;
signal \DFT.done_c_0\ : std_logic;
signal \DFT.o_done_RNOZ0Z_0_cascade_\ : std_logic;
signal done_c : std_logic;
signal \INVDFT.o_doneC_net\ : std_logic;
signal \DFT.state_RNIHM3GZ0Z_0\ : std_logic;
signal \o_X_c_18\ : std_logic;
signal \o_X_c_16\ : std_logic;
signal \INVo_X_1__nesr_2C_net\ : std_logic;
signal \o_X_c_19\ : std_logic;
signal \INVo_X_1__nesr_3C_net\ : std_logic;
signal \o_X_c_21\ : std_logic;
signal \INVo_X_1__nesr_5C_net\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_2\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_2\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_619\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_1\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_620\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_1\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_621\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_0\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_622\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_ma_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_4\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_4\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_625\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_626\ : std_logic;
signal \bfn_9_20_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_627\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_628\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO\ : std_logic;
signal \X_1__8\ : std_logic;
signal \INVDFT.o_X_1__nesr_8C_net\ : std_logic;
signal \X_1__9\ : std_logic;
signal \INVDFT.o_X_1__nesr_7C_net\ : std_logic;
signal \X_1__7\ : std_logic;
signal \o_X_c_17\ : std_logic;
signal \o_X_c_23\ : std_logic;
signal \INVo_X_1__nesr_1C_net\ : std_logic;
signal \bfn_10_17_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_583\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_584\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_585\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_586\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_ma_1\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_5\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_5\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_589\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_590\ : std_logic;
signal \bfn_10_18_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_591\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_592\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_593\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_594\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_2\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_3\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_2\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_583_THRU_CO\ : std_logic;
signal \bfn_10_19_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_584_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_4\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_585_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_3_3\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_586_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_2\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_587\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_3\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_588\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_6_1\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_589_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_7_1\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_590_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_8_1\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_9_0\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_591_THRU_CO\ : std_logic;
signal \bfn_10_20_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_592_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_10_0\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_593_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_11\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_axb_9\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_12\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_621_THRU_CO\ : std_logic;
signal \bfn_10_21_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_622_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_3\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_623\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_3_2\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_624\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_1\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_625_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_2\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_626_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_6_0\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_627_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_7_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_8\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_8_THRU_CO\ : std_logic;
signal \X_1__6\ : std_logic;
signal \bfn_10_22_0_\ : std_logic;
signal \INVDFT.o_X_1__nesr_6C_net\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_620_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_824\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_1\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNI8J5C1\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_825\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_3_0\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_826\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_860\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_8\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_827\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_861\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_1\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_828\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_862\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_6\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_829\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_863\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_7\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_830\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_864\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_8_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_9\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_831\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_865\ : std_logic;
signal \bfn_10_23_0_\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_axb_11\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_10\ : std_logic;
signal \X_1__11\ : std_logic;
signal \X_1__13\ : std_logic;
signal \INVDFT.o_X_1__nesr_12C_net\ : std_logic;
signal \X_1__12\ : std_logic;
signal \o_X_c_22\ : std_logic;
signal \INVo_X_1__nesr_6C_net\ : std_logic;
signal \o_X_c_20\ : std_logic;
signal \INVo_X_1__nesr_4C_net\ : std_logic;
signal \bfn_11_17_0_\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_1\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_549_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_549\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_550_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_550\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_551\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_6\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_552\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_6\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_553_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_553\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_554\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_554_THRU_CO\ : std_logic;
signal \bfn_11_18_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_555_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_555\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_556_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_556\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_557_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_557\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_558_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_558\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_559_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_559\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_594_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_560\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_axb_13\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_3\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_655_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_655\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_656_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_656\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_657_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_657\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_658_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_658\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_659\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_7\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_660\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_7\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_661_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_661\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_662\ : std_logic;
signal \bfn_11_20_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_662_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_13_0_c_RNO\ : std_logic;
signal \DFT.state_2_0_cascade_\ : std_logic;
signal \INVDFT.state_0C_net\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO\ : std_logic;
signal \DFT.x_7\ : std_logic;
signal \DFT.x_9\ : std_logic;
signal \DFT.x_8\ : std_logic;
signal \INVDFT.o_X_0__nesr_7C_net\ : std_logic;
signal \bfn_11_22_0_\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_THRU_CO\ : std_logic;
signal \X_1__10\ : std_logic;
signal \bfn_11_23_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_964\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_0\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_965\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_3\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_966\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNIRG904\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_967\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_axb_7\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_6_2\ : std_logic;
signal \INVDFT.o_X_1__nesr_10C_net\ : std_logic;
signal \DFT.un1_state_1_0\ : std_logic;
signal \DFT.x_13\ : std_logic;
signal \DFT.x_12\ : std_logic;
signal \DFT.x_15\ : std_logic;
signal \INVDFT.o_X_0__nesr_13C_net\ : std_logic;
signal \X_0__15\ : std_logic;
signal \o_X_c_15\ : std_logic;
signal \INVo_X_0__nesr_9C_net\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_3\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_3\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_4\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_4\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_1\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_6_b_l_ofx\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_6_ma_1\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_2\ : std_logic;
signal \DFT.stateZ0Z_0\ : std_logic;
signal i_rst_c : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_1\ : std_logic;
signal \DFT.state_2_0\ : std_logic;
signal \DFT.stateZ0Z_1\ : std_logic;
signal \INVDFT.b_6C_net\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_1\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_1\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_ma_2\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_5_b_l_ofx_2\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_6_ma_2\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_5\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_4\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_ma_3\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_4\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_3\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_5\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_763_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_763\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_764\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_axb_3\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_963\ : std_logic;
signal \INVDFT.o_X_0__nesr_10C_net\ : std_logic;
signal \DFT.x_14\ : std_logic;
signal \INVDFT.o_X_0__nesr_14C_net\ : std_logic;
signal \DFT.x_11\ : std_logic;
signal \INVDFT.o_X_0__nesr_11C_net\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_897\ : std_logic;
signal \bfn_13_17_0_\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_898\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_2\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_899\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_3_1\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_6_a\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_900\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_5_b_l_ofx_1\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_6_ma_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_12_0_c_RNO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_2\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_5_b_l_ofx_0\ : std_logic;
signal \DFT.bZ0Z_6\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_6_ma\ : std_logic;
signal \DFT.aZ0Z_0\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_0\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_823\ : std_logic;
signal \INVDFT.o_X_0__nesr_6C_net\ : std_logic;
signal \DFT.un1_state_4_0\ : std_logic;
signal \X_0__13\ : std_logic;
signal \o_X_c_7\ : std_logic;
signal \INVo_X_0__nesr_7C_net\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_0\ : std_logic;
signal \bfn_14_17_0_\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_0\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_727_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_727\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_728_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_728\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_729_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_729\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_730\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_730_THRU_CO\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_1\ : std_logic;
signal \bfn_14_18_0_\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_1\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_691\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_0\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_692_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_692\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_0\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_693\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_694_THRU_CO\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_694\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_5_b_l_ofx\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_ma\ : std_logic;
signal \DFT.multiplier.mult1_AdderTree2i_bigtree_695\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_4_3\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5\ : std_logic;
signal \DFT.multiplier.regsA_un3_result_cry_5_THRU_CO\ : std_logic;
signal \X_0__7\ : std_logic;
signal \o_X_c_1\ : std_logic;
signal \X_0__6\ : std_logic;
signal \o_X_c_0\ : std_logic;
signal \INVo_X_0__nesr_1C_net\ : std_logic;
signal \X_1__14\ : std_logic;
signal \o_X_c_24\ : std_logic;
signal \INVo_X_1__nesr_8C_net\ : std_logic;
signal \X_0__9\ : std_logic;
signal \o_X_c_3\ : std_logic;
signal \X_0__8\ : std_logic;
signal \o_X_c_2\ : std_logic;
signal \INVo_X_0__nesr_3C_net\ : std_logic;
signal \X_0__10\ : std_logic;
signal \o_X_c_4\ : std_logic;
signal \INVo_X_0__nesr_4C_net\ : std_logic;
signal \X_0__14\ : std_logic;
signal \o_X_c_8\ : std_logic;
signal \INVo_X_0__nesr_8C_net\ : std_logic;
signal \X_1__15\ : std_logic;
signal \o_X_c_31\ : std_logic;
signal \INVo_X_1__nesr_9C_net\ : std_logic;
signal \X_0__11\ : std_logic;
signal \o_X_c_5\ : std_logic;
signal \X_0__12\ : std_logic;
signal \o_X_c_6\ : std_logic;
signal \INVo_X_0__nesr_5C_net\ : std_logic;
signal done_c_0_g : std_logic;
signal i_rst_c_i_g : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \o_X_wire\ : std_logic_vector(31 downto 0);
signal i_ref_clk_wire : std_logic;
signal i_rst_wire : std_logic;
signal done_wire : std_logic;
signal \pll_DYNAMICDELAY_wire\ : std_logic_vector(7 downto 0);

begin
    o_X <= \o_X_wire\;
    i_ref_clk_wire <= i_ref_clk;
    i_rst_wire <= i_rst;
    done <= done_wire;
    \pll_DYNAMICDELAY_wire\ <= \GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\&\GNDG0\;

    \pll\ : SB_PLL40_CORE
    generic map (
            DELAY_ADJUSTMENT_MODE_FEEDBACK => "FIXED",
            TEST_MODE => '0',
            SHIFTREG_DIV_MODE => "00",
            PLLOUT_SELECT => "GENCLK",
            FILTER_RANGE => "010",
            FEEDBACK_PATH => "SIMPLE",
            FDA_RELATIVE => "0000",
            FDA_FEEDBACK => "0000",
            ENABLE_ICEGATE => '0',
            DIVR => "0100",
            DIVQ => "101",
            DIVF => "0101111",
            DELAY_ADJUSTMENT_MODE_RELATIVE => "FIXED"
        )
    port map (
            EXTFEEDBACK => '0',
            LATCHINPUTVALUE => '0',
            SCLK => '0',
            SDO => OPEN,
            LOCK => OPEN,
            PLLOUTCORE => sys_clk,
            REFERENCECLK => \N__3401\,
            RESETB => \N__6419\,
            BYPASS => \GNDG0\,
            SDI => '0',
            DYNAMICDELAY => \pll_DYNAMICDELAY_wire\,
            PLLOUTGLOBAL => OPEN
        );

    \o_X_obuf_29_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7068\,
            DIN => \N__7067\,
            DOUT => \N__7066\,
            PACKAGEPIN => \o_X_wire\(29)
        );

    \o_X_obuf_29_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7068\,
            PADOUT => \N__7067\,
            PADIN => \N__7066\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6695\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_9_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7059\,
            DIN => \N__7058\,
            DOUT => \N__7057\,
            PACKAGEPIN => \o_X_wire\(9)
        );

    \o_X_obuf_9_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7059\,
            PADOUT => \N__7058\,
            PADIN => \N__7057\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4968\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_26_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7050\,
            DIN => \N__7049\,
            DOUT => \N__7048\,
            PACKAGEPIN => \o_X_wire\(26)
        );

    \o_X_obuf_26_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7050\,
            PADOUT => \N__7049\,
            PADIN => \N__7048\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6684\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_ref_clk_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7041\,
            DIN => \N__7040\,
            DOUT => \N__7039\,
            PACKAGEPIN => i_ref_clk_wire
        );

    \i_ref_clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__7041\,
            PADOUT => \N__7040\,
            PADIN => \N__7039\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_ref_clk_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_31_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7032\,
            DIN => \N__7031\,
            DOUT => \N__7030\,
            PACKAGEPIN => \o_X_wire\(31)
        );

    \o_X_obuf_31_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7032\,
            PADOUT => \N__7031\,
            PADIN => \N__7030\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6697\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7023\,
            DIN => \N__7022\,
            DOUT => \N__7021\,
            PACKAGEPIN => \o_X_wire\(7)
        );

    \o_X_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7023\,
            PADOUT => \N__7022\,
            PADIN => \N__7021\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__5570\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_13_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7014\,
            DIN => \N__7013\,
            DOUT => \N__7012\,
            PACKAGEPIN => \o_X_wire\(13)
        );

    \o_X_obuf_13_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7014\,
            PADOUT => \N__7013\,
            PADIN => \N__7012\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4938\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__7005\,
            DIN => \N__7004\,
            DOUT => \N__7003\,
            PACKAGEPIN => \o_X_wire\(2)
        );

    \o_X_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__7005\,
            PADOUT => \N__7004\,
            PADIN => \N__7003\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6248\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_14_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6996\,
            DIN => \N__6995\,
            DOUT => \N__6994\,
            PACKAGEPIN => \o_X_wire\(14)
        );

    \o_X_obuf_14_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6996\,
            PADOUT => \N__6995\,
            PADIN => \N__6994\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4958\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_24_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6987\,
            DIN => \N__6986\,
            DOUT => \N__6985\,
            PACKAGEPIN => \o_X_wire\(24)
        );

    \o_X_obuf_24_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6987\,
            PADOUT => \N__6986\,
            PADIN => \N__6985\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6299\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \i_rst_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6978\,
            DIN => \N__6977\,
            DOUT => \N__6976\,
            PACKAGEPIN => i_rst_wire
        );

    \i_rst_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__6978\,
            PADOUT => \N__6977\,
            PADIN => \N__6976\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => i_rst_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6969\,
            DIN => \N__6968\,
            DOUT => \N__6967\,
            PACKAGEPIN => \o_X_wire\(5)
        );

    \o_X_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6969\,
            PADOUT => \N__6968\,
            PADIN => \N__6967\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6620\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_11_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6960\,
            DIN => \N__6959\,
            DOUT => \N__6958\,
            PACKAGEPIN => \o_X_wire\(11)
        );

    \o_X_obuf_11_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6960\,
            PADOUT => \N__6959\,
            PADIN => \N__6958\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4975\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_27_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6951\,
            DIN => \N__6950\,
            DOUT => \N__6949\,
            PACKAGEPIN => \o_X_wire\(27)
        );

    \o_X_obuf_27_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6951\,
            PADOUT => \N__6950\,
            PADIN => \N__6949\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6683\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_0_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6942\,
            DIN => \N__6941\,
            DOUT => \N__6940\,
            PACKAGEPIN => \o_X_wire\(0)
        );

    \o_X_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6942\,
            PADOUT => \N__6941\,
            PADIN => \N__6940\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6332\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_22_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6933\,
            DIN => \N__6932\,
            DOUT => \N__6931\,
            PACKAGEPIN => \o_X_wire\(22)
        );

    \o_X_obuf_22_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6933\,
            PADOUT => \N__6932\,
            PADIN => \N__6931\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4274\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_19_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6924\,
            DIN => \N__6923\,
            DOUT => \N__6922\,
            PACKAGEPIN => \o_X_wire\(19)
        );

    \o_X_obuf_19_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6924\,
            PADOUT => \N__6923\,
            PADIN => \N__6922\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3434\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_28_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6915\,
            DIN => \N__6914\,
            DOUT => \N__6913\,
            PACKAGEPIN => \o_X_wire\(28)
        );

    \o_X_obuf_28_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6915\,
            PADOUT => \N__6914\,
            PADIN => \N__6913\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6696\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_30_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6906\,
            DIN => \N__6905\,
            DOUT => \N__6904\,
            PACKAGEPIN => \o_X_wire\(30)
        );

    \o_X_obuf_30_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6906\,
            PADOUT => \N__6905\,
            PADIN => \N__6904\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6698\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_8_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6897\,
            DIN => \N__6896\,
            DOUT => \N__6895\,
            PACKAGEPIN => \o_X_wire\(8)
        );

    \o_X_obuf_8_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6897\,
            PADOUT => \N__6896\,
            PADIN => \N__6895\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6731\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \done_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6888\,
            DIN => \N__6887\,
            DOUT => \N__6886\,
            PACKAGEPIN => done_wire
        );

    \done_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6888\,
            PADOUT => \N__6887\,
            PADIN => \N__6886\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3527\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_12_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6879\,
            DIN => \N__6878\,
            DOUT => \N__6877\,
            PACKAGEPIN => \o_X_wire\(12)
        );

    \o_X_obuf_12_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6879\,
            PADOUT => \N__6878\,
            PADIN => \N__6877\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4959\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6870\,
            DIN => \N__6869\,
            DOUT => \N__6868\,
            PACKAGEPIN => \o_X_wire\(3)
        );

    \o_X_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6870\,
            PADOUT => \N__6869\,
            PADIN => \N__6868\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6269\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_17_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6861\,
            DIN => \N__6860\,
            DOUT => \N__6859\,
            PACKAGEPIN => \o_X_wire\(17)
        );

    \o_X_obuf_17_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6861\,
            PADOUT => \N__6860\,
            PADIN => \N__6859\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3677\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_25_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6852\,
            DIN => \N__6851\,
            DOUT => \N__6850\,
            PACKAGEPIN => \o_X_wire\(25)
        );

    \o_X_obuf_25_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6852\,
            PADOUT => \N__6851\,
            PADIN => \N__6850\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6685\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_20_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6843\,
            DIN => \N__6842\,
            DOUT => \N__6841\,
            PACKAGEPIN => \o_X_wire\(20)
        );

    \o_X_obuf_20_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6843\,
            PADOUT => \N__6842\,
            PADIN => \N__6841\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4262\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6834\,
            DIN => \N__6833\,
            DOUT => \N__6832\,
            PACKAGEPIN => \o_X_wire\(6)
        );

    \o_X_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6834\,
            PADOUT => \N__6833\,
            PADIN => \N__6832\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6596\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_10_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6825\,
            DIN => \N__6824\,
            DOUT => \N__6823\,
            PACKAGEPIN => \o_X_wire\(10)
        );

    \o_X_obuf_10_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6825\,
            PADOUT => \N__6824\,
            PADIN => \N__6823\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4976\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6816\,
            DIN => \N__6815\,
            DOUT => \N__6814\,
            PACKAGEPIN => \o_X_wire\(1)
        );

    \o_X_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6816\,
            PADOUT => \N__6815\,
            PADIN => \N__6814\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6359\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_15_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6807\,
            DIN => \N__6806\,
            DOUT => \N__6805\,
            PACKAGEPIN => \o_X_wire\(15)
        );

    \o_X_obuf_15_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6807\,
            PADOUT => \N__6806\,
            PADIN => \N__6805\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__4937\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_23_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6798\,
            DIN => \N__6797\,
            DOUT => \N__6796\,
            PACKAGEPIN => \o_X_wire\(23)
        );

    \o_X_obuf_23_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6798\,
            PADOUT => \N__6797\,
            PADIN => \N__6796\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3659\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_18_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6789\,
            DIN => \N__6788\,
            DOUT => \N__6787\,
            PACKAGEPIN => \o_X_wire\(18)
        );

    \o_X_obuf_18_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6789\,
            PADOUT => \N__6788\,
            PADIN => \N__6787\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3470\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6780\,
            DIN => \N__6779\,
            DOUT => \N__6778\,
            PACKAGEPIN => \o_X_wire\(4)
        );

    \o_X_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6780\,
            PADOUT => \N__6779\,
            PADIN => \N__6778\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6224\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_16_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6771\,
            DIN => \N__6770\,
            DOUT => \N__6769\,
            PACKAGEPIN => \o_X_wire\(16)
        );

    \o_X_obuf_16_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6771\,
            PADOUT => \N__6770\,
            PADIN => \N__6769\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3452\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \o_X_obuf_21_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__6762\,
            DIN => \N__6761\,
            DOUT => \N__6760\,
            PACKAGEPIN => \o_X_wire\(21)
        );

    \o_X_obuf_21_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__6762\,
            PADOUT => \N__6761\,
            PADIN => \N__6760\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3419\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__1467\ : InMux
    port map (
            O => \N__6743\,
            I => \N__6740\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__6740\,
            I => \N__6737\
        );

    \I__1465\ : Span4Mux_h
    port map (
            O => \N__6737\,
            I => \N__6734\
        );

    \I__1464\ : Odrv4
    port map (
            O => \N__6734\,
            I => \X_0__14\
        );

    \I__1463\ : IoInMux
    port map (
            O => \N__6731\,
            I => \N__6728\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6728\,
            I => \N__6725\
        );

    \I__1461\ : Span4Mux_s0_v
    port map (
            O => \N__6725\,
            I => \N__6722\
        );

    \I__1460\ : Span4Mux_h
    port map (
            O => \N__6722\,
            I => \N__6719\
        );

    \I__1459\ : Span4Mux_v
    port map (
            O => \N__6719\,
            I => \N__6716\
        );

    \I__1458\ : Span4Mux_v
    port map (
            O => \N__6716\,
            I => \N__6713\
        );

    \I__1457\ : Odrv4
    port map (
            O => \N__6713\,
            I => \o_X_c_8\
        );

    \I__1456\ : InMux
    port map (
            O => \N__6710\,
            I => \N__6707\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__6707\,
            I => \N__6704\
        );

    \I__1454\ : Span4Mux_h
    port map (
            O => \N__6704\,
            I => \N__6701\
        );

    \I__1453\ : Odrv4
    port map (
            O => \N__6701\,
            I => \X_1__15\
        );

    \I__1452\ : IoInMux
    port map (
            O => \N__6698\,
            I => \N__6692\
        );

    \I__1451\ : IoInMux
    port map (
            O => \N__6697\,
            I => \N__6689\
        );

    \I__1450\ : IoInMux
    port map (
            O => \N__6696\,
            I => \N__6686\
        );

    \I__1449\ : IoInMux
    port map (
            O => \N__6695\,
            I => \N__6680\
        );

    \I__1448\ : LocalMux
    port map (
            O => \N__6692\,
            I => \N__6673\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__6689\,
            I => \N__6673\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__6686\,
            I => \N__6673\
        );

    \I__1445\ : IoInMux
    port map (
            O => \N__6685\,
            I => \N__6670\
        );

    \I__1444\ : IoInMux
    port map (
            O => \N__6684\,
            I => \N__6667\
        );

    \I__1443\ : IoInMux
    port map (
            O => \N__6683\,
            I => \N__6664\
        );

    \I__1442\ : LocalMux
    port map (
            O => \N__6680\,
            I => \N__6661\
        );

    \I__1441\ : IoSpan4Mux
    port map (
            O => \N__6673\,
            I => \N__6652\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__6670\,
            I => \N__6652\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6667\,
            I => \N__6652\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__6664\,
            I => \N__6652\
        );

    \I__1437\ : Span4Mux_s3_h
    port map (
            O => \N__6661\,
            I => \N__6649\
        );

    \I__1436\ : IoSpan4Mux
    port map (
            O => \N__6652\,
            I => \N__6646\
        );

    \I__1435\ : Span4Mux_v
    port map (
            O => \N__6649\,
            I => \N__6641\
        );

    \I__1434\ : Span4Mux_s3_h
    port map (
            O => \N__6646\,
            I => \N__6641\
        );

    \I__1433\ : Sp12to4
    port map (
            O => \N__6641\,
            I => \N__6638\
        );

    \I__1432\ : Span12Mux_h
    port map (
            O => \N__6638\,
            I => \N__6635\
        );

    \I__1431\ : Span12Mux_v
    port map (
            O => \N__6635\,
            I => \N__6632\
        );

    \I__1430\ : Odrv12
    port map (
            O => \N__6632\,
            I => \o_X_c_31\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6629\,
            I => \N__6626\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__6626\,
            I => \N__6623\
        );

    \I__1427\ : Odrv12
    port map (
            O => \N__6623\,
            I => \X_0__11\
        );

    \I__1426\ : IoInMux
    port map (
            O => \N__6620\,
            I => \N__6617\
        );

    \I__1425\ : LocalMux
    port map (
            O => \N__6617\,
            I => \N__6614\
        );

    \I__1424\ : Sp12to4
    port map (
            O => \N__6614\,
            I => \N__6611\
        );

    \I__1423\ : Span12Mux_h
    port map (
            O => \N__6611\,
            I => \N__6608\
        );

    \I__1422\ : Odrv12
    port map (
            O => \N__6608\,
            I => \o_X_c_5\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6605\,
            I => \N__6602\
        );

    \I__1420\ : LocalMux
    port map (
            O => \N__6602\,
            I => \N__6599\
        );

    \I__1419\ : Odrv12
    port map (
            O => \N__6599\,
            I => \X_0__12\
        );

    \I__1418\ : IoInMux
    port map (
            O => \N__6596\,
            I => \N__6593\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6593\,
            I => \N__6590\
        );

    \I__1416\ : Span12Mux_s5_h
    port map (
            O => \N__6590\,
            I => \N__6587\
        );

    \I__1415\ : Span12Mux_h
    port map (
            O => \N__6587\,
            I => \N__6584\
        );

    \I__1414\ : Odrv12
    port map (
            O => \N__6584\,
            I => \o_X_c_6\
        );

    \I__1413\ : CEMux
    port map (
            O => \N__6581\,
            I => \N__6536\
        );

    \I__1412\ : CEMux
    port map (
            O => \N__6580\,
            I => \N__6536\
        );

    \I__1411\ : CEMux
    port map (
            O => \N__6579\,
            I => \N__6536\
        );

    \I__1410\ : CEMux
    port map (
            O => \N__6578\,
            I => \N__6536\
        );

    \I__1409\ : CEMux
    port map (
            O => \N__6577\,
            I => \N__6536\
        );

    \I__1408\ : CEMux
    port map (
            O => \N__6576\,
            I => \N__6536\
        );

    \I__1407\ : CEMux
    port map (
            O => \N__6575\,
            I => \N__6536\
        );

    \I__1406\ : CEMux
    port map (
            O => \N__6574\,
            I => \N__6536\
        );

    \I__1405\ : CEMux
    port map (
            O => \N__6573\,
            I => \N__6536\
        );

    \I__1404\ : CEMux
    port map (
            O => \N__6572\,
            I => \N__6536\
        );

    \I__1403\ : CEMux
    port map (
            O => \N__6571\,
            I => \N__6536\
        );

    \I__1402\ : CEMux
    port map (
            O => \N__6570\,
            I => \N__6536\
        );

    \I__1401\ : CEMux
    port map (
            O => \N__6569\,
            I => \N__6536\
        );

    \I__1400\ : CEMux
    port map (
            O => \N__6568\,
            I => \N__6536\
        );

    \I__1399\ : CEMux
    port map (
            O => \N__6567\,
            I => \N__6536\
        );

    \I__1398\ : GlobalMux
    port map (
            O => \N__6536\,
            I => \N__6533\
        );

    \I__1397\ : gio2CtrlBuf
    port map (
            O => \N__6533\,
            I => done_c_0_g
        );

    \I__1396\ : InMux
    port map (
            O => \N__6530\,
            I => \N__6525\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6529\,
            I => \N__6522\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6528\,
            I => \N__6519\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__6525\,
            I => \N__6492\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__6522\,
            I => \N__6487\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__6519\,
            I => \N__6484\
        );

    \I__1390\ : SRMux
    port map (
            O => \N__6518\,
            I => \N__6425\
        );

    \I__1389\ : SRMux
    port map (
            O => \N__6517\,
            I => \N__6425\
        );

    \I__1388\ : SRMux
    port map (
            O => \N__6516\,
            I => \N__6425\
        );

    \I__1387\ : SRMux
    port map (
            O => \N__6515\,
            I => \N__6425\
        );

    \I__1386\ : SRMux
    port map (
            O => \N__6514\,
            I => \N__6425\
        );

    \I__1385\ : SRMux
    port map (
            O => \N__6513\,
            I => \N__6425\
        );

    \I__1384\ : SRMux
    port map (
            O => \N__6512\,
            I => \N__6425\
        );

    \I__1383\ : SRMux
    port map (
            O => \N__6511\,
            I => \N__6425\
        );

    \I__1382\ : SRMux
    port map (
            O => \N__6510\,
            I => \N__6425\
        );

    \I__1381\ : SRMux
    port map (
            O => \N__6509\,
            I => \N__6425\
        );

    \I__1380\ : SRMux
    port map (
            O => \N__6508\,
            I => \N__6425\
        );

    \I__1379\ : SRMux
    port map (
            O => \N__6507\,
            I => \N__6425\
        );

    \I__1378\ : SRMux
    port map (
            O => \N__6506\,
            I => \N__6425\
        );

    \I__1377\ : SRMux
    port map (
            O => \N__6505\,
            I => \N__6425\
        );

    \I__1376\ : SRMux
    port map (
            O => \N__6504\,
            I => \N__6425\
        );

    \I__1375\ : SRMux
    port map (
            O => \N__6503\,
            I => \N__6425\
        );

    \I__1374\ : SRMux
    port map (
            O => \N__6502\,
            I => \N__6425\
        );

    \I__1373\ : SRMux
    port map (
            O => \N__6501\,
            I => \N__6425\
        );

    \I__1372\ : SRMux
    port map (
            O => \N__6500\,
            I => \N__6425\
        );

    \I__1371\ : SRMux
    port map (
            O => \N__6499\,
            I => \N__6425\
        );

    \I__1370\ : SRMux
    port map (
            O => \N__6498\,
            I => \N__6425\
        );

    \I__1369\ : SRMux
    port map (
            O => \N__6497\,
            I => \N__6425\
        );

    \I__1368\ : SRMux
    port map (
            O => \N__6496\,
            I => \N__6425\
        );

    \I__1367\ : SRMux
    port map (
            O => \N__6495\,
            I => \N__6425\
        );

    \I__1366\ : Glb2LocalMux
    port map (
            O => \N__6492\,
            I => \N__6425\
        );

    \I__1365\ : SRMux
    port map (
            O => \N__6491\,
            I => \N__6425\
        );

    \I__1364\ : SRMux
    port map (
            O => \N__6490\,
            I => \N__6425\
        );

    \I__1363\ : Glb2LocalMux
    port map (
            O => \N__6487\,
            I => \N__6425\
        );

    \I__1362\ : Glb2LocalMux
    port map (
            O => \N__6484\,
            I => \N__6425\
        );

    \I__1361\ : GlobalMux
    port map (
            O => \N__6425\,
            I => \N__6422\
        );

    \I__1360\ : gio2CtrlBuf
    port map (
            O => \N__6422\,
            I => i_rst_c_i_g
        );

    \I__1359\ : IoInMux
    port map (
            O => \N__6419\,
            I => \N__6416\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__6416\,
            I => \N__6413\
        );

    \I__1357\ : IoSpan4Mux
    port map (
            O => \N__6413\,
            I => \N__6410\
        );

    \I__1356\ : Span4Mux_s0_v
    port map (
            O => \N__6410\,
            I => \N__6407\
        );

    \I__1355\ : Odrv4
    port map (
            O => \N__6407\,
            I => \CONSTANT_ONE_NET\
        );

    \I__1354\ : InMux
    port map (
            O => \N__6404\,
            I => \N__6401\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__6401\,
            I => \DFT.multiplier.regsA_un3_result_5_b_l_ofx\
        );

    \I__1352\ : CascadeMux
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6395\,
            I => \N__6392\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6392\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_ma\
        );

    \I__1349\ : InMux
    port map (
            O => \N__6389\,
            I => \N__6386\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__6386\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_695\
        );

    \I__1347\ : InMux
    port map (
            O => \N__6383\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_3\
        );

    \I__1346\ : InMux
    port map (
            O => \N__6380\,
            I => \DFT.multiplier.regsA_un3_result_cry_5\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6377\,
            I => \N__6374\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6374\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_THRU_CO\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6371\,
            I => \N__6368\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6368\,
            I => \N__6365\
        );

    \I__1341\ : Span4Mux_h
    port map (
            O => \N__6365\,
            I => \N__6362\
        );

    \I__1340\ : Odrv4
    port map (
            O => \N__6362\,
            I => \X_0__7\
        );

    \I__1339\ : IoInMux
    port map (
            O => \N__6359\,
            I => \N__6356\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6356\,
            I => \N__6353\
        );

    \I__1337\ : IoSpan4Mux
    port map (
            O => \N__6353\,
            I => \N__6350\
        );

    \I__1336\ : Span4Mux_s1_h
    port map (
            O => \N__6350\,
            I => \N__6347\
        );

    \I__1335\ : Sp12to4
    port map (
            O => \N__6347\,
            I => \N__6344\
        );

    \I__1334\ : Span12Mux_h
    port map (
            O => \N__6344\,
            I => \N__6341\
        );

    \I__1333\ : Odrv12
    port map (
            O => \N__6341\,
            I => \o_X_c_1\
        );

    \I__1332\ : InMux
    port map (
            O => \N__6338\,
            I => \N__6335\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__6335\,
            I => \X_0__6\
        );

    \I__1330\ : IoInMux
    port map (
            O => \N__6332\,
            I => \N__6329\
        );

    \I__1329\ : LocalMux
    port map (
            O => \N__6329\,
            I => \N__6326\
        );

    \I__1328\ : Span4Mux_s2_h
    port map (
            O => \N__6326\,
            I => \N__6323\
        );

    \I__1327\ : Span4Mux_h
    port map (
            O => \N__6323\,
            I => \N__6320\
        );

    \I__1326\ : Sp12to4
    port map (
            O => \N__6320\,
            I => \N__6317\
        );

    \I__1325\ : Span12Mux_v
    port map (
            O => \N__6317\,
            I => \N__6314\
        );

    \I__1324\ : Odrv12
    port map (
            O => \N__6314\,
            I => \o_X_c_0\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6308\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6308\,
            I => \N__6305\
        );

    \I__1321\ : Span4Mux_h
    port map (
            O => \N__6305\,
            I => \N__6302\
        );

    \I__1320\ : Odrv4
    port map (
            O => \N__6302\,
            I => \X_1__14\
        );

    \I__1319\ : IoInMux
    port map (
            O => \N__6299\,
            I => \N__6296\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6296\,
            I => \N__6293\
        );

    \I__1317\ : Span4Mux_s2_h
    port map (
            O => \N__6293\,
            I => \N__6290\
        );

    \I__1316\ : Sp12to4
    port map (
            O => \N__6290\,
            I => \N__6287\
        );

    \I__1315\ : Span12Mux_v
    port map (
            O => \N__6287\,
            I => \N__6284\
        );

    \I__1314\ : Span12Mux_h
    port map (
            O => \N__6284\,
            I => \N__6281\
        );

    \I__1313\ : Odrv12
    port map (
            O => \N__6281\,
            I => \o_X_c_24\
        );

    \I__1312\ : InMux
    port map (
            O => \N__6278\,
            I => \N__6275\
        );

    \I__1311\ : LocalMux
    port map (
            O => \N__6275\,
            I => \N__6272\
        );

    \I__1310\ : Odrv4
    port map (
            O => \N__6272\,
            I => \X_0__9\
        );

    \I__1309\ : IoInMux
    port map (
            O => \N__6269\,
            I => \N__6266\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6266\,
            I => \N__6263\
        );

    \I__1307\ : Span12Mux_s10_h
    port map (
            O => \N__6263\,
            I => \N__6260\
        );

    \I__1306\ : Odrv12
    port map (
            O => \N__6260\,
            I => \o_X_c_3\
        );

    \I__1305\ : InMux
    port map (
            O => \N__6257\,
            I => \N__6254\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__6254\,
            I => \N__6251\
        );

    \I__1303\ : Odrv4
    port map (
            O => \N__6251\,
            I => \X_0__8\
        );

    \I__1302\ : IoInMux
    port map (
            O => \N__6248\,
            I => \N__6245\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__6245\,
            I => \N__6242\
        );

    \I__1300\ : Span12Mux_s9_h
    port map (
            O => \N__6242\,
            I => \N__6239\
        );

    \I__1299\ : Odrv12
    port map (
            O => \N__6239\,
            I => \o_X_c_2\
        );

    \I__1298\ : InMux
    port map (
            O => \N__6236\,
            I => \N__6233\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__6233\,
            I => \N__6230\
        );

    \I__1296\ : Span4Mux_h
    port map (
            O => \N__6230\,
            I => \N__6227\
        );

    \I__1295\ : Odrv4
    port map (
            O => \N__6227\,
            I => \X_0__10\
        );

    \I__1294\ : IoInMux
    port map (
            O => \N__6224\,
            I => \N__6221\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6221\,
            I => \N__6218\
        );

    \I__1292\ : Span12Mux_s10_h
    port map (
            O => \N__6218\,
            I => \N__6215\
        );

    \I__1291\ : Odrv12
    port map (
            O => \N__6215\,
            I => \o_X_c_4\
        );

    \I__1290\ : InMux
    port map (
            O => \N__6212\,
            I => \N__6209\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6209\,
            I => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO\
        );

    \I__1288\ : CascadeMux
    port map (
            O => \N__6206\,
            I => \N__6203\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6203\,
            I => \N__6200\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6200\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_728_THRU_CO\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6197\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_728\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6191\
        );

    \I__1283\ : LocalMux
    port map (
            O => \N__6191\,
            I => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__6188\,
            I => \N__6185\
        );

    \I__1281\ : InMux
    port map (
            O => \N__6185\,
            I => \N__6182\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__6182\,
            I => \N__6179\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__6179\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_729_THRU_CO\
        );

    \I__1278\ : InMux
    port map (
            O => \N__6176\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_729\
        );

    \I__1277\ : InMux
    port map (
            O => \N__6173\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_730\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6167\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__6167\,
            I => \N__6164\
        );

    \I__1274\ : Odrv4
    port map (
            O => \N__6164\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_730_THRU_CO\
        );

    \I__1273\ : CascadeMux
    port map (
            O => \N__6161\,
            I => \N__6158\
        );

    \I__1272\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6155\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__6155\,
            I => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_1\
        );

    \I__1270\ : CascadeMux
    port map (
            O => \N__6152\,
            I => \N__6149\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6149\,
            I => \N__6146\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6146\,
            I => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_1\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6143\,
            I => \N__6139\
        );

    \I__1266\ : InMux
    port map (
            O => \N__6142\,
            I => \N__6136\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6139\,
            I => \N__6133\
        );

    \I__1264\ : LocalMux
    port map (
            O => \N__6136\,
            I => \N__6130\
        );

    \I__1263\ : Span4Mux_h
    port map (
            O => \N__6133\,
            I => \N__6127\
        );

    \I__1262\ : Span4Mux_v
    port map (
            O => \N__6130\,
            I => \N__6124\
        );

    \I__1261\ : Span4Mux_v
    port map (
            O => \N__6127\,
            I => \N__6121\
        );

    \I__1260\ : Odrv4
    port map (
            O => \N__6124\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_CO\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__6121\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_CO\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6116\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_691\
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__6113\,
            I => \N__6110\
        );

    \I__1256\ : InMux
    port map (
            O => \N__6110\,
            I => \N__6107\
        );

    \I__1255\ : LocalMux
    port map (
            O => \N__6107\,
            I => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_0\
        );

    \I__1254\ : InMux
    port map (
            O => \N__6104\,
            I => \N__6101\
        );

    \I__1253\ : LocalMux
    port map (
            O => \N__6101\,
            I => \N__6098\
        );

    \I__1252\ : Span4Mux_v
    port map (
            O => \N__6098\,
            I => \N__6095\
        );

    \I__1251\ : Span4Mux_h
    port map (
            O => \N__6095\,
            I => \N__6092\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__6092\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_692_THRU_CO\
        );

    \I__1249\ : InMux
    port map (
            O => \N__6089\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_692\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__6086\,
            I => \N__6083\
        );

    \I__1247\ : InMux
    port map (
            O => \N__6083\,
            I => \N__6080\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__6080\,
            I => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_0\
        );

    \I__1245\ : CascadeMux
    port map (
            O => \N__6077\,
            I => \N__6073\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6076\,
            I => \N__6070\
        );

    \I__1243\ : InMux
    port map (
            O => \N__6073\,
            I => \N__6067\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__6070\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_CO\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6067\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_CO\
        );

    \I__1240\ : InMux
    port map (
            O => \N__6062\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_693\
        );

    \I__1239\ : InMux
    port map (
            O => \N__6059\,
            I => \N__6056\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__6056\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO\
        );

    \I__1237\ : InMux
    port map (
            O => \N__6053\,
            I => \N__6050\
        );

    \I__1236\ : LocalMux
    port map (
            O => \N__6050\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_694_THRU_CO\
        );

    \I__1235\ : InMux
    port map (
            O => \N__6047\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_694\
        );

    \I__1234\ : InMux
    port map (
            O => \N__6044\,
            I => \N__6041\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__6041\,
            I => \N__6038\
        );

    \I__1232\ : Odrv12
    port map (
            O => \N__6038\,
            I => \DFT.multiplier.regsA_un3_result_5_b_l_ofx_0\
        );

    \I__1231\ : InMux
    port map (
            O => \N__6035\,
            I => \N__6029\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__6034\,
            I => \N__6023\
        );

    \I__1229\ : CascadeMux
    port map (
            O => \N__6033\,
            I => \N__6019\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__6032\,
            I => \N__6015\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__6029\,
            I => \N__6010\
        );

    \I__1226\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6007\
        );

    \I__1225\ : InMux
    port map (
            O => \N__6027\,
            I => \N__6002\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6026\,
            I => \N__6002\
        );

    \I__1223\ : InMux
    port map (
            O => \N__6023\,
            I => \N__5997\
        );

    \I__1222\ : InMux
    port map (
            O => \N__6022\,
            I => \N__5997\
        );

    \I__1221\ : InMux
    port map (
            O => \N__6019\,
            I => \N__5992\
        );

    \I__1220\ : InMux
    port map (
            O => \N__6018\,
            I => \N__5992\
        );

    \I__1219\ : InMux
    port map (
            O => \N__6015\,
            I => \N__5989\
        );

    \I__1218\ : InMux
    port map (
            O => \N__6014\,
            I => \N__5984\
        );

    \I__1217\ : InMux
    port map (
            O => \N__6013\,
            I => \N__5984\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__6010\,
            I => \DFT.bZ0Z_6\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__6007\,
            I => \DFT.bZ0Z_6\
        );

    \I__1214\ : LocalMux
    port map (
            O => \N__6002\,
            I => \DFT.bZ0Z_6\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__5997\,
            I => \DFT.bZ0Z_6\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5992\,
            I => \DFT.bZ0Z_6\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5989\,
            I => \DFT.bZ0Z_6\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__5984\,
            I => \DFT.bZ0Z_6\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__5969\,
            I => \N__5966\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5966\,
            I => \N__5963\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__5963\,
            I => \N__5960\
        );

    \I__1206\ : Span4Mux_h
    port map (
            O => \N__5960\,
            I => \N__5957\
        );

    \I__1205\ : Odrv4
    port map (
            O => \N__5957\,
            I => \DFT.multiplier.regsA_un3_result_cry_6_ma\
        );

    \I__1204\ : CascadeMux
    port map (
            O => \N__5954\,
            I => \N__5948\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5953\,
            I => \N__5936\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5952\,
            I => \N__5936\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5951\,
            I => \N__5922\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5913\
        );

    \I__1199\ : InMux
    port map (
            O => \N__5947\,
            I => \N__5913\
        );

    \I__1198\ : InMux
    port map (
            O => \N__5946\,
            I => \N__5913\
        );

    \I__1197\ : InMux
    port map (
            O => \N__5945\,
            I => \N__5913\
        );

    \I__1196\ : InMux
    port map (
            O => \N__5944\,
            I => \N__5908\
        );

    \I__1195\ : InMux
    port map (
            O => \N__5943\,
            I => \N__5908\
        );

    \I__1194\ : InMux
    port map (
            O => \N__5942\,
            I => \N__5903\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5941\,
            I => \N__5903\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5936\,
            I => \N__5865\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5935\,
            I => \N__5848\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5934\,
            I => \N__5848\
        );

    \I__1189\ : InMux
    port map (
            O => \N__5933\,
            I => \N__5848\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5932\,
            I => \N__5848\
        );

    \I__1187\ : InMux
    port map (
            O => \N__5931\,
            I => \N__5848\
        );

    \I__1186\ : InMux
    port map (
            O => \N__5930\,
            I => \N__5848\
        );

    \I__1185\ : InMux
    port map (
            O => \N__5929\,
            I => \N__5848\
        );

    \I__1184\ : InMux
    port map (
            O => \N__5928\,
            I => \N__5848\
        );

    \I__1183\ : InMux
    port map (
            O => \N__5927\,
            I => \N__5841\
        );

    \I__1182\ : InMux
    port map (
            O => \N__5926\,
            I => \N__5841\
        );

    \I__1181\ : InMux
    port map (
            O => \N__5925\,
            I => \N__5841\
        );

    \I__1180\ : LocalMux
    port map (
            O => \N__5922\,
            I => \N__5826\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__5913\,
            I => \N__5826\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5908\,
            I => \N__5826\
        );

    \I__1177\ : LocalMux
    port map (
            O => \N__5903\,
            I => \N__5823\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5902\,
            I => \N__5808\
        );

    \I__1175\ : InMux
    port map (
            O => \N__5901\,
            I => \N__5808\
        );

    \I__1174\ : InMux
    port map (
            O => \N__5900\,
            I => \N__5808\
        );

    \I__1173\ : InMux
    port map (
            O => \N__5899\,
            I => \N__5808\
        );

    \I__1172\ : InMux
    port map (
            O => \N__5898\,
            I => \N__5808\
        );

    \I__1171\ : InMux
    port map (
            O => \N__5897\,
            I => \N__5808\
        );

    \I__1170\ : InMux
    port map (
            O => \N__5896\,
            I => \N__5808\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5895\,
            I => \N__5791\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5894\,
            I => \N__5791\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5893\,
            I => \N__5791\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5892\,
            I => \N__5791\
        );

    \I__1165\ : InMux
    port map (
            O => \N__5891\,
            I => \N__5791\
        );

    \I__1164\ : InMux
    port map (
            O => \N__5890\,
            I => \N__5791\
        );

    \I__1163\ : InMux
    port map (
            O => \N__5889\,
            I => \N__5791\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5888\,
            I => \N__5791\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5887\,
            I => \N__5774\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5886\,
            I => \N__5774\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5885\,
            I => \N__5774\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5884\,
            I => \N__5774\
        );

    \I__1157\ : InMux
    port map (
            O => \N__5883\,
            I => \N__5774\
        );

    \I__1156\ : InMux
    port map (
            O => \N__5882\,
            I => \N__5774\
        );

    \I__1155\ : InMux
    port map (
            O => \N__5881\,
            I => \N__5774\
        );

    \I__1154\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5774\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5759\
        );

    \I__1152\ : InMux
    port map (
            O => \N__5878\,
            I => \N__5759\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5759\
        );

    \I__1150\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5759\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5759\
        );

    \I__1148\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5759\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5873\,
            I => \N__5759\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5872\,
            I => \N__5750\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5871\,
            I => \N__5750\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5870\,
            I => \N__5750\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5869\,
            I => \N__5750\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5868\,
            I => \N__5747\
        );

    \I__1141\ : Span4Mux_v
    port map (
            O => \N__5865\,
            I => \N__5740\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5848\,
            I => \N__5740\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5841\,
            I => \N__5740\
        );

    \I__1138\ : InMux
    port map (
            O => \N__5840\,
            I => \N__5723\
        );

    \I__1137\ : InMux
    port map (
            O => \N__5839\,
            I => \N__5723\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5838\,
            I => \N__5723\
        );

    \I__1135\ : InMux
    port map (
            O => \N__5837\,
            I => \N__5723\
        );

    \I__1134\ : InMux
    port map (
            O => \N__5836\,
            I => \N__5723\
        );

    \I__1133\ : InMux
    port map (
            O => \N__5835\,
            I => \N__5723\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5834\,
            I => \N__5723\
        );

    \I__1131\ : InMux
    port map (
            O => \N__5833\,
            I => \N__5723\
        );

    \I__1130\ : Odrv4
    port map (
            O => \N__5826\,
            I => \DFT.aZ0Z_0\
        );

    \I__1129\ : Odrv4
    port map (
            O => \N__5823\,
            I => \DFT.aZ0Z_0\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__5808\,
            I => \DFT.aZ0Z_0\
        );

    \I__1127\ : LocalMux
    port map (
            O => \N__5791\,
            I => \DFT.aZ0Z_0\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5774\,
            I => \DFT.aZ0Z_0\
        );

    \I__1125\ : LocalMux
    port map (
            O => \N__5759\,
            I => \DFT.aZ0Z_0\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5750\,
            I => \DFT.aZ0Z_0\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__5747\,
            I => \DFT.aZ0Z_0\
        );

    \I__1122\ : Odrv4
    port map (
            O => \N__5740\,
            I => \DFT.aZ0Z_0\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__5723\,
            I => \DFT.aZ0Z_0\
        );

    \I__1120\ : CascadeMux
    port map (
            O => \N__5702\,
            I => \N__5699\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5699\,
            I => \N__5696\
        );

    \I__1118\ : LocalMux
    port map (
            O => \N__5696\,
            I => \N__5693\
        );

    \I__1117\ : Span4Mux_h
    port map (
            O => \N__5693\,
            I => \N__5690\
        );

    \I__1116\ : Odrv4
    port map (
            O => \N__5690\,
            I => \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_0\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5687\,
            I => \N__5683\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5686\,
            I => \N__5680\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5683\,
            I => \N__5677\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__5680\,
            I => \N__5674\
        );

    \I__1111\ : Span4Mux_h
    port map (
            O => \N__5677\,
            I => \N__5671\
        );

    \I__1110\ : Span4Mux_v
    port map (
            O => \N__5674\,
            I => \N__5668\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__5671\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_CO\
        );

    \I__1108\ : Odrv4
    port map (
            O => \N__5668\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_CO\
        );

    \I__1107\ : InMux
    port map (
            O => \N__5663\,
            I => \N__5659\
        );

    \I__1106\ : CascadeMux
    port map (
            O => \N__5662\,
            I => \N__5656\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5659\,
            I => \N__5653\
        );

    \I__1104\ : InMux
    port map (
            O => \N__5656\,
            I => \N__5650\
        );

    \I__1103\ : Span4Mux_h
    port map (
            O => \N__5653\,
            I => \N__5647\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__5650\,
            I => \N__5644\
        );

    \I__1101\ : Odrv4
    port map (
            O => \N__5647\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_823\
        );

    \I__1100\ : Odrv4
    port map (
            O => \N__5644\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_823\
        );

    \I__1099\ : CEMux
    port map (
            O => \N__5639\,
            I => \N__5635\
        );

    \I__1098\ : CEMux
    port map (
            O => \N__5638\,
            I => \N__5629\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5635\,
            I => \N__5626\
        );

    \I__1096\ : CEMux
    port map (
            O => \N__5634\,
            I => \N__5623\
        );

    \I__1095\ : CEMux
    port map (
            O => \N__5633\,
            I => \N__5619\
        );

    \I__1094\ : CEMux
    port map (
            O => \N__5632\,
            I => \N__5616\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__5629\,
            I => \N__5609\
        );

    \I__1092\ : Span4Mux_h
    port map (
            O => \N__5626\,
            I => \N__5609\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5623\,
            I => \N__5609\
        );

    \I__1090\ : CEMux
    port map (
            O => \N__5622\,
            I => \N__5606\
        );

    \I__1089\ : LocalMux
    port map (
            O => \N__5619\,
            I => \N__5601\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__5616\,
            I => \N__5601\
        );

    \I__1087\ : Span4Mux_v
    port map (
            O => \N__5609\,
            I => \N__5596\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5606\,
            I => \N__5596\
        );

    \I__1085\ : Span4Mux_v
    port map (
            O => \N__5601\,
            I => \N__5593\
        );

    \I__1084\ : Span4Mux_h
    port map (
            O => \N__5596\,
            I => \N__5590\
        );

    \I__1083\ : Span4Mux_h
    port map (
            O => \N__5593\,
            I => \N__5587\
        );

    \I__1082\ : Odrv4
    port map (
            O => \N__5590\,
            I => \DFT.un1_state_4_0\
        );

    \I__1081\ : Odrv4
    port map (
            O => \N__5587\,
            I => \DFT.un1_state_4_0\
        );

    \I__1080\ : InMux
    port map (
            O => \N__5582\,
            I => \N__5579\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5579\,
            I => \N__5576\
        );

    \I__1078\ : Span4Mux_v
    port map (
            O => \N__5576\,
            I => \N__5573\
        );

    \I__1077\ : Odrv4
    port map (
            O => \N__5573\,
            I => \X_0__13\
        );

    \I__1076\ : IoInMux
    port map (
            O => \N__5570\,
            I => \N__5567\
        );

    \I__1075\ : LocalMux
    port map (
            O => \N__5567\,
            I => \N__5564\
        );

    \I__1074\ : Span4Mux_s2_v
    port map (
            O => \N__5564\,
            I => \N__5561\
        );

    \I__1073\ : Span4Mux_v
    port map (
            O => \N__5561\,
            I => \N__5558\
        );

    \I__1072\ : Sp12to4
    port map (
            O => \N__5558\,
            I => \N__5555\
        );

    \I__1071\ : Span12Mux_s9_h
    port map (
            O => \N__5555\,
            I => \N__5552\
        );

    \I__1070\ : Odrv12
    port map (
            O => \N__5552\,
            I => \o_X_c_7\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__5549\,
            I => \N__5546\
        );

    \I__1068\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5543\
        );

    \I__1067\ : LocalMux
    port map (
            O => \N__5543\,
            I => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_0\
        );

    \I__1066\ : CascadeMux
    port map (
            O => \N__5540\,
            I => \N__5537\
        );

    \I__1065\ : InMux
    port map (
            O => \N__5537\,
            I => \N__5534\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__5534\,
            I => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_0\
        );

    \I__1063\ : InMux
    port map (
            O => \N__5531\,
            I => \N__5528\
        );

    \I__1062\ : LocalMux
    port map (
            O => \N__5528\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_727_THRU_CO\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5525\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_727\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5522\,
            I => \N__5519\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5519\,
            I => \N__5516\
        );

    \I__1058\ : Span4Mux_v
    port map (
            O => \N__5516\,
            I => \N__5513\
        );

    \I__1057\ : Odrv4
    port map (
            O => \N__5513\,
            I => \DFT.multiplier.regsA_un3_result_cry_12_0_c_RNO\
        );

    \I__1056\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5507\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5507\,
            I => \N__5504\
        );

    \I__1054\ : Span4Mux_h
    port map (
            O => \N__5504\,
            I => \N__5501\
        );

    \I__1053\ : Odrv4
    port map (
            O => \N__5501\,
            I => \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_0\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5495\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5495\,
            I => \N__5492\
        );

    \I__1050\ : Odrv4
    port map (
            O => \N__5492\,
            I => \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_2\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5489\,
            I => \N__5486\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5486\,
            I => \N__5483\
        );

    \I__1047\ : Span4Mux_h
    port map (
            O => \N__5483\,
            I => \N__5480\
        );

    \I__1046\ : Span4Mux_v
    port map (
            O => \N__5480\,
            I => \N__5477\
        );

    \I__1045\ : Odrv4
    port map (
            O => \N__5477\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_897\
        );

    \I__1044\ : InMux
    port map (
            O => \N__5474\,
            I => \N__5471\
        );

    \I__1043\ : LocalMux
    port map (
            O => \N__5471\,
            I => \N__5468\
        );

    \I__1042\ : Span4Mux_h
    port map (
            O => \N__5468\,
            I => \N__5465\
        );

    \I__1041\ : Span4Mux_v
    port map (
            O => \N__5465\,
            I => \N__5462\
        );

    \I__1040\ : Odrv4
    port map (
            O => \N__5462\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_898\
        );

    \I__1039\ : InMux
    port map (
            O => \N__5459\,
            I => \DFT.multiplier.regsA_un3_result_cry_2_2\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__5456\,
            I => \N__5453\
        );

    \I__1037\ : InMux
    port map (
            O => \N__5453\,
            I => \N__5450\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5450\,
            I => \N__5447\
        );

    \I__1035\ : Span4Mux_h
    port map (
            O => \N__5447\,
            I => \N__5444\
        );

    \I__1034\ : Span4Mux_v
    port map (
            O => \N__5444\,
            I => \N__5441\
        );

    \I__1033\ : Odrv4
    port map (
            O => \N__5441\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_899\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5438\,
            I => \DFT.multiplier.regsA_un3_result_cry_3_1\
        );

    \I__1031\ : CascadeMux
    port map (
            O => \N__5435\,
            I => \N__5432\
        );

    \I__1030\ : InMux
    port map (
            O => \N__5432\,
            I => \N__5429\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5429\,
            I => \DFT.multiplier.regsA_un3_result_6_a\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5426\,
            I => \DFT.multiplier.regsA_un3_result_cry_4\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5423\,
            I => \N__5420\
        );

    \I__1026\ : LocalMux
    port map (
            O => \N__5420\,
            I => \N__5417\
        );

    \I__1025\ : Odrv4
    port map (
            O => \N__5417\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_900\
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__5414\,
            I => \N__5411\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5411\,
            I => \N__5408\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__5408\,
            I => \N__5405\
        );

    \I__1021\ : Odrv4
    port map (
            O => \N__5405\,
            I => \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_0\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5402\,
            I => \N__5399\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5399\,
            I => \N__5396\
        );

    \I__1018\ : Odrv4
    port map (
            O => \N__5396\,
            I => \DFT.multiplier.regsA_un3_result_5_b_l_ofx_1\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__5393\,
            I => \N__5390\
        );

    \I__1016\ : InMux
    port map (
            O => \N__5390\,
            I => \N__5387\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5387\,
            I => \N__5384\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__5384\,
            I => \DFT.multiplier.regsA_un3_result_cry_6_ma_0\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5381\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_764\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5378\,
            I => \N__5375\
        );

    \I__1011\ : LocalMux
    port map (
            O => \N__5375\,
            I => \N__5372\
        );

    \I__1010\ : Span4Mux_h
    port map (
            O => \N__5372\,
            I => \N__5369\
        );

    \I__1009\ : Odrv4
    port map (
            O => \N__5369\,
            I => \DFT.multiplier.regsA_un3_result_axb_3\
        );

    \I__1008\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5363\
        );

    \I__1007\ : LocalMux
    port map (
            O => \N__5363\,
            I => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__5360\,
            I => \N__5357\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5354\
        );

    \I__1004\ : LocalMux
    port map (
            O => \N__5354\,
            I => \N__5351\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__5351\,
            I => \DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO_0\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5348\,
            I => \N__5345\
        );

    \I__1001\ : LocalMux
    port map (
            O => \N__5345\,
            I => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5338\
        );

    \I__999\ : CascadeMux
    port map (
            O => \N__5341\,
            I => \N__5335\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__5338\,
            I => \N__5332\
        );

    \I__997\ : InMux
    port map (
            O => \N__5335\,
            I => \N__5329\
        );

    \I__996\ : Odrv4
    port map (
            O => \N__5332\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_963\
        );

    \I__995\ : LocalMux
    port map (
            O => \N__5329\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_963\
        );

    \I__994\ : InMux
    port map (
            O => \N__5324\,
            I => \N__5320\
        );

    \I__993\ : InMux
    port map (
            O => \N__5323\,
            I => \N__5317\
        );

    \I__992\ : LocalMux
    port map (
            O => \N__5320\,
            I => \DFT.x_14\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5317\,
            I => \DFT.x_14\
        );

    \I__990\ : CascadeMux
    port map (
            O => \N__5312\,
            I => \N__5309\
        );

    \I__989\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5305\
        );

    \I__988\ : InMux
    port map (
            O => \N__5308\,
            I => \N__5302\
        );

    \I__987\ : LocalMux
    port map (
            O => \N__5305\,
            I => \DFT.x_11\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__5302\,
            I => \DFT.x_11\
        );

    \I__985\ : InMux
    port map (
            O => \N__5297\,
            I => \N__5294\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5294\,
            I => \DFT.multiplier.regsA_un3_result_cry_6_ma_2\
        );

    \I__983\ : CascadeMux
    port map (
            O => \N__5291\,
            I => \N__5288\
        );

    \I__982\ : InMux
    port map (
            O => \N__5288\,
            I => \N__5285\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5285\,
            I => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_5\
        );

    \I__980\ : CascadeMux
    port map (
            O => \N__5282\,
            I => \N__5279\
        );

    \I__979\ : InMux
    port map (
            O => \N__5279\,
            I => \N__5276\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5276\,
            I => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_4\
        );

    \I__977\ : CascadeMux
    port map (
            O => \N__5273\,
            I => \N__5270\
        );

    \I__976\ : InMux
    port map (
            O => \N__5270\,
            I => \N__5267\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__5267\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_ma_3\
        );

    \I__974\ : CascadeMux
    port map (
            O => \N__5264\,
            I => \N__5261\
        );

    \I__973\ : InMux
    port map (
            O => \N__5261\,
            I => \N__5258\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__5258\,
            I => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_4\
        );

    \I__971\ : CascadeMux
    port map (
            O => \N__5255\,
            I => \N__5252\
        );

    \I__970\ : InMux
    port map (
            O => \N__5252\,
            I => \N__5249\
        );

    \I__969\ : LocalMux
    port map (
            O => \N__5249\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_3\
        );

    \I__968\ : CascadeMux
    port map (
            O => \N__5246\,
            I => \N__5243\
        );

    \I__967\ : InMux
    port map (
            O => \N__5243\,
            I => \N__5240\
        );

    \I__966\ : LocalMux
    port map (
            O => \N__5240\,
            I => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_5\
        );

    \I__965\ : InMux
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__5234\,
            I => \N__5231\
        );

    \I__963\ : Span4Mux_h
    port map (
            O => \N__5231\,
            I => \N__5228\
        );

    \I__962\ : Odrv4
    port map (
            O => \N__5228\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_763_THRU_CO\
        );

    \I__961\ : InMux
    port map (
            O => \N__5225\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_763\
        );

    \I__960\ : InMux
    port map (
            O => \N__5222\,
            I => \N__5218\
        );

    \I__959\ : InMux
    port map (
            O => \N__5221\,
            I => \N__5214\
        );

    \I__958\ : LocalMux
    port map (
            O => \N__5218\,
            I => \N__5211\
        );

    \I__957\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5208\
        );

    \I__956\ : LocalMux
    port map (
            O => \N__5214\,
            I => \N__5204\
        );

    \I__955\ : Span4Mux_h
    port map (
            O => \N__5211\,
            I => \N__5201\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__5208\,
            I => \N__5198\
        );

    \I__953\ : InMux
    port map (
            O => \N__5207\,
            I => \N__5195\
        );

    \I__952\ : Odrv4
    port map (
            O => \N__5204\,
            I => \DFT.stateZ0Z_0\
        );

    \I__951\ : Odrv4
    port map (
            O => \N__5201\,
            I => \DFT.stateZ0Z_0\
        );

    \I__950\ : Odrv12
    port map (
            O => \N__5198\,
            I => \DFT.stateZ0Z_0\
        );

    \I__949\ : LocalMux
    port map (
            O => \N__5195\,
            I => \DFT.stateZ0Z_0\
        );

    \I__948\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5183\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__5183\,
            I => \N__5180\
        );

    \I__946\ : Span4Mux_v
    port map (
            O => \N__5180\,
            I => \N__5175\
        );

    \I__945\ : InMux
    port map (
            O => \N__5179\,
            I => \N__5172\
        );

    \I__944\ : InMux
    port map (
            O => \N__5178\,
            I => \N__5168\
        );

    \I__943\ : Span4Mux_h
    port map (
            O => \N__5175\,
            I => \N__5160\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5172\,
            I => \N__5160\
        );

    \I__941\ : CascadeMux
    port map (
            O => \N__5171\,
            I => \N__5157\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5168\,
            I => \N__5154\
        );

    \I__939\ : InMux
    port map (
            O => \N__5167\,
            I => \N__5147\
        );

    \I__938\ : InMux
    port map (
            O => \N__5166\,
            I => \N__5147\
        );

    \I__937\ : InMux
    port map (
            O => \N__5165\,
            I => \N__5147\
        );

    \I__936\ : Span4Mux_h
    port map (
            O => \N__5160\,
            I => \N__5144\
        );

    \I__935\ : InMux
    port map (
            O => \N__5157\,
            I => \N__5141\
        );

    \I__934\ : Span4Mux_v
    port map (
            O => \N__5154\,
            I => \N__5138\
        );

    \I__933\ : LocalMux
    port map (
            O => \N__5147\,
            I => \N__5135\
        );

    \I__932\ : Span4Mux_h
    port map (
            O => \N__5144\,
            I => \N__5130\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__5141\,
            I => \N__5130\
        );

    \I__930\ : Span4Mux_h
    port map (
            O => \N__5138\,
            I => \N__5125\
        );

    \I__929\ : Span4Mux_v
    port map (
            O => \N__5135\,
            I => \N__5125\
        );

    \I__928\ : Span4Mux_v
    port map (
            O => \N__5130\,
            I => \N__5122\
        );

    \I__927\ : Sp12to4
    port map (
            O => \N__5125\,
            I => \N__5119\
        );

    \I__926\ : Span4Mux_h
    port map (
            O => \N__5122\,
            I => \N__5116\
        );

    \I__925\ : Span12Mux_h
    port map (
            O => \N__5119\,
            I => \N__5111\
        );

    \I__924\ : Sp12to4
    port map (
            O => \N__5116\,
            I => \N__5111\
        );

    \I__923\ : Span12Mux_v
    port map (
            O => \N__5111\,
            I => \N__5108\
        );

    \I__922\ : Odrv12
    port map (
            O => \N__5108\,
            I => i_rst_c
        );

    \I__921\ : CascadeMux
    port map (
            O => \N__5105\,
            I => \N__5102\
        );

    \I__920\ : InMux
    port map (
            O => \N__5102\,
            I => \N__5099\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__5099\,
            I => \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_1\
        );

    \I__918\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__917\ : LocalMux
    port map (
            O => \N__5093\,
            I => \N__5088\
        );

    \I__916\ : InMux
    port map (
            O => \N__5092\,
            I => \N__5083\
        );

    \I__915\ : InMux
    port map (
            O => \N__5091\,
            I => \N__5083\
        );

    \I__914\ : Odrv4
    port map (
            O => \N__5088\,
            I => \DFT.state_2_0\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5083\,
            I => \DFT.state_2_0\
        );

    \I__912\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5073\
        );

    \I__911\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5067\
        );

    \I__910\ : InMux
    port map (
            O => \N__5076\,
            I => \N__5067\
        );

    \I__909\ : LocalMux
    port map (
            O => \N__5073\,
            I => \N__5062\
        );

    \I__908\ : InMux
    port map (
            O => \N__5072\,
            I => \N__5059\
        );

    \I__907\ : LocalMux
    port map (
            O => \N__5067\,
            I => \N__5056\
        );

    \I__906\ : InMux
    port map (
            O => \N__5066\,
            I => \N__5051\
        );

    \I__905\ : InMux
    port map (
            O => \N__5065\,
            I => \N__5051\
        );

    \I__904\ : Span4Mux_h
    port map (
            O => \N__5062\,
            I => \N__5048\
        );

    \I__903\ : LocalMux
    port map (
            O => \N__5059\,
            I => \N__5045\
        );

    \I__902\ : Odrv4
    port map (
            O => \N__5056\,
            I => \DFT.stateZ0Z_1\
        );

    \I__901\ : LocalMux
    port map (
            O => \N__5051\,
            I => \DFT.stateZ0Z_1\
        );

    \I__900\ : Odrv4
    port map (
            O => \N__5048\,
            I => \DFT.stateZ0Z_1\
        );

    \I__899\ : Odrv12
    port map (
            O => \N__5045\,
            I => \DFT.stateZ0Z_1\
        );

    \I__898\ : CascadeMux
    port map (
            O => \N__5036\,
            I => \N__5033\
        );

    \I__897\ : InMux
    port map (
            O => \N__5033\,
            I => \N__5030\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__5030\,
            I => \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_1\
        );

    \I__895\ : CascadeMux
    port map (
            O => \N__5027\,
            I => \N__5024\
        );

    \I__894\ : InMux
    port map (
            O => \N__5024\,
            I => \N__5021\
        );

    \I__893\ : LocalMux
    port map (
            O => \N__5021\,
            I => \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_1\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__5018\,
            I => \N__5015\
        );

    \I__891\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5012\
        );

    \I__890\ : LocalMux
    port map (
            O => \N__5012\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_ma_2\
        );

    \I__889\ : CascadeMux
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__888\ : InMux
    port map (
            O => \N__5006\,
            I => \N__5003\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5003\,
            I => \DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO_0\
        );

    \I__886\ : InMux
    port map (
            O => \N__5000\,
            I => \N__4997\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4997\,
            I => \N__4994\
        );

    \I__884\ : Odrv4
    port map (
            O => \N__4994\,
            I => \DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO\
        );

    \I__883\ : InMux
    port map (
            O => \N__4991\,
            I => \N__4988\
        );

    \I__882\ : LocalMux
    port map (
            O => \N__4988\,
            I => \DFT.multiplier.regsA_un3_result_5_b_l_ofx_2\
        );

    \I__881\ : InMux
    port map (
            O => \N__4985\,
            I => \N__4982\
        );

    \I__880\ : LocalMux
    port map (
            O => \N__4982\,
            I => \N__4979\
        );

    \I__879\ : Odrv4
    port map (
            O => \N__4979\,
            I => \X_0__15\
        );

    \I__878\ : IoInMux
    port map (
            O => \N__4976\,
            I => \N__4972\
        );

    \I__877\ : IoInMux
    port map (
            O => \N__4975\,
            I => \N__4969\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__4972\,
            I => \N__4963\
        );

    \I__875\ : LocalMux
    port map (
            O => \N__4969\,
            I => \N__4963\
        );

    \I__874\ : IoInMux
    port map (
            O => \N__4968\,
            I => \N__4960\
        );

    \I__873\ : IoSpan4Mux
    port map (
            O => \N__4963\,
            I => \N__4955\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4960\,
            I => \N__4952\
        );

    \I__871\ : IoInMux
    port map (
            O => \N__4959\,
            I => \N__4949\
        );

    \I__870\ : IoInMux
    port map (
            O => \N__4958\,
            I => \N__4946\
        );

    \I__869\ : IoSpan4Mux
    port map (
            O => \N__4955\,
            I => \N__4939\
        );

    \I__868\ : IoSpan4Mux
    port map (
            O => \N__4952\,
            I => \N__4939\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4949\,
            I => \N__4939\
        );

    \I__866\ : LocalMux
    port map (
            O => \N__4946\,
            I => \N__4934\
        );

    \I__865\ : IoSpan4Mux
    port map (
            O => \N__4939\,
            I => \N__4931\
        );

    \I__864\ : IoInMux
    port map (
            O => \N__4938\,
            I => \N__4928\
        );

    \I__863\ : IoInMux
    port map (
            O => \N__4937\,
            I => \N__4925\
        );

    \I__862\ : IoSpan4Mux
    port map (
            O => \N__4934\,
            I => \N__4922\
        );

    \I__861\ : Span4Mux_s3_v
    port map (
            O => \N__4931\,
            I => \N__4919\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4928\,
            I => \N__4916\
        );

    \I__859\ : LocalMux
    port map (
            O => \N__4925\,
            I => \N__4913\
        );

    \I__858\ : IoSpan4Mux
    port map (
            O => \N__4922\,
            I => \N__4910\
        );

    \I__857\ : Span4Mux_v
    port map (
            O => \N__4919\,
            I => \N__4905\
        );

    \I__856\ : Span4Mux_s3_v
    port map (
            O => \N__4916\,
            I => \N__4905\
        );

    \I__855\ : Span12Mux_s6_v
    port map (
            O => \N__4913\,
            I => \N__4902\
        );

    \I__854\ : Span4Mux_s3_v
    port map (
            O => \N__4910\,
            I => \N__4897\
        );

    \I__853\ : Span4Mux_h
    port map (
            O => \N__4905\,
            I => \N__4897\
        );

    \I__852\ : Odrv12
    port map (
            O => \N__4902\,
            I => \o_X_c_15\
        );

    \I__851\ : Odrv4
    port map (
            O => \N__4897\,
            I => \o_X_c_15\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__4892\,
            I => \N__4889\
        );

    \I__849\ : InMux
    port map (
            O => \N__4889\,
            I => \N__4886\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4886\,
            I => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_3\
        );

    \I__847\ : CascadeMux
    port map (
            O => \N__4883\,
            I => \N__4880\
        );

    \I__846\ : InMux
    port map (
            O => \N__4880\,
            I => \N__4877\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4877\,
            I => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_3\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__4874\,
            I => \N__4871\
        );

    \I__843\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4868\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4868\,
            I => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_4\
        );

    \I__841\ : CascadeMux
    port map (
            O => \N__4865\,
            I => \N__4862\
        );

    \I__840\ : InMux
    port map (
            O => \N__4862\,
            I => \N__4859\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__4859\,
            I => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_4\
        );

    \I__838\ : CascadeMux
    port map (
            O => \N__4856\,
            I => \N__4853\
        );

    \I__837\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4850\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4850\,
            I => \N__4847\
        );

    \I__835\ : Odrv4
    port map (
            O => \N__4847\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_1\
        );

    \I__834\ : CascadeMux
    port map (
            O => \N__4844\,
            I => \N__4841\
        );

    \I__833\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4838\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4838\,
            I => \DFT.multiplier.regsA_un3_result_6_b_l_ofx\
        );

    \I__831\ : InMux
    port map (
            O => \N__4835\,
            I => \N__4832\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4832\,
            I => \DFT.multiplier.regsA_un3_result_cry_6_ma_1\
        );

    \I__829\ : CascadeMux
    port map (
            O => \N__4829\,
            I => \N__4826\
        );

    \I__828\ : InMux
    port map (
            O => \N__4826\,
            I => \N__4823\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4823\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_2\
        );

    \I__826\ : CascadeMux
    port map (
            O => \N__4820\,
            I => \N__4817\
        );

    \I__825\ : InMux
    port map (
            O => \N__4817\,
            I => \N__4814\
        );

    \I__824\ : LocalMux
    port map (
            O => \N__4814\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_965\
        );

    \I__823\ : InMux
    port map (
            O => \N__4811\,
            I => \DFT.multiplier.regsA_un3_result_cry_3\
        );

    \I__822\ : CascadeMux
    port map (
            O => \N__4808\,
            I => \N__4805\
        );

    \I__821\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4802\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4802\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_966\
        );

    \I__819\ : InMux
    port map (
            O => \N__4799\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_0\
        );

    \I__818\ : InMux
    port map (
            O => \N__4796\,
            I => \N__4793\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4793\,
            I => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNIRG904\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__4790\,
            I => \N__4786\
        );

    \I__815\ : InMux
    port map (
            O => \N__4789\,
            I => \N__4783\
        );

    \I__814\ : InMux
    port map (
            O => \N__4786\,
            I => \N__4780\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4783\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_967\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__4780\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_967\
        );

    \I__811\ : InMux
    port map (
            O => \N__4775\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_0\
        );

    \I__810\ : InMux
    port map (
            O => \N__4772\,
            I => \N__4769\
        );

    \I__809\ : LocalMux
    port map (
            O => \N__4769\,
            I => \DFT.multiplier.regsA_un3_result_axb_7\
        );

    \I__808\ : InMux
    port map (
            O => \N__4766\,
            I => \DFT.multiplier.regsA_un3_result_cry_6_2\
        );

    \I__807\ : CEMux
    port map (
            O => \N__4763\,
            I => \N__4759\
        );

    \I__806\ : CEMux
    port map (
            O => \N__4762\,
            I => \N__4755\
        );

    \I__805\ : LocalMux
    port map (
            O => \N__4759\,
            I => \N__4752\
        );

    \I__804\ : CEMux
    port map (
            O => \N__4758\,
            I => \N__4747\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4755\,
            I => \N__4744\
        );

    \I__802\ : Span4Mux_v
    port map (
            O => \N__4752\,
            I => \N__4741\
        );

    \I__801\ : CEMux
    port map (
            O => \N__4751\,
            I => \N__4738\
        );

    \I__800\ : CEMux
    port map (
            O => \N__4750\,
            I => \N__4735\
        );

    \I__799\ : LocalMux
    port map (
            O => \N__4747\,
            I => \N__4732\
        );

    \I__798\ : Span4Mux_v
    port map (
            O => \N__4744\,
            I => \N__4725\
        );

    \I__797\ : Span4Mux_h
    port map (
            O => \N__4741\,
            I => \N__4725\
        );

    \I__796\ : LocalMux
    port map (
            O => \N__4738\,
            I => \N__4725\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__4735\,
            I => \N__4722\
        );

    \I__794\ : Span4Mux_h
    port map (
            O => \N__4732\,
            I => \N__4719\
        );

    \I__793\ : Span4Mux_h
    port map (
            O => \N__4725\,
            I => \N__4716\
        );

    \I__792\ : Span4Mux_h
    port map (
            O => \N__4722\,
            I => \N__4713\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__4719\,
            I => \DFT.un1_state_1_0\
        );

    \I__790\ : Odrv4
    port map (
            O => \N__4716\,
            I => \DFT.un1_state_1_0\
        );

    \I__789\ : Odrv4
    port map (
            O => \N__4713\,
            I => \DFT.un1_state_1_0\
        );

    \I__788\ : InMux
    port map (
            O => \N__4706\,
            I => \N__4702\
        );

    \I__787\ : InMux
    port map (
            O => \N__4705\,
            I => \N__4699\
        );

    \I__786\ : LocalMux
    port map (
            O => \N__4702\,
            I => \DFT.x_13\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4699\,
            I => \DFT.x_13\
        );

    \I__784\ : InMux
    port map (
            O => \N__4694\,
            I => \N__4690\
        );

    \I__783\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4687\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4690\,
            I => \DFT.x_12\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4687\,
            I => \DFT.x_12\
        );

    \I__780\ : InMux
    port map (
            O => \N__4682\,
            I => \N__4678\
        );

    \I__779\ : InMux
    port map (
            O => \N__4681\,
            I => \N__4675\
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4678\,
            I => \DFT.x_15\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4675\,
            I => \DFT.x_15\
        );

    \I__776\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4667\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4667\,
            I => \N__4664\
        );

    \I__774\ : Span4Mux_h
    port map (
            O => \N__4664\,
            I => \N__4661\
        );

    \I__773\ : Odrv4
    port map (
            O => \N__4661\,
            I => \DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO\
        );

    \I__772\ : InMux
    port map (
            O => \N__4658\,
            I => \N__4654\
        );

    \I__771\ : InMux
    port map (
            O => \N__4657\,
            I => \N__4651\
        );

    \I__770\ : LocalMux
    port map (
            O => \N__4654\,
            I => \DFT.x_7\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4651\,
            I => \DFT.x_7\
        );

    \I__768\ : InMux
    port map (
            O => \N__4646\,
            I => \N__4642\
        );

    \I__767\ : InMux
    port map (
            O => \N__4645\,
            I => \N__4639\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4642\,
            I => \DFT.x_9\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4639\,
            I => \DFT.x_9\
        );

    \I__764\ : InMux
    port map (
            O => \N__4634\,
            I => \N__4630\
        );

    \I__763\ : InMux
    port map (
            O => \N__4633\,
            I => \N__4627\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4630\,
            I => \DFT.x_8\
        );

    \I__761\ : LocalMux
    port map (
            O => \N__4627\,
            I => \DFT.x_8\
        );

    \I__760\ : InMux
    port map (
            O => \N__4622\,
            I => \DFT.multiplier.regsA_un3_result_cry_2\
        );

    \I__759\ : CascadeMux
    port map (
            O => \N__4619\,
            I => \N__4616\
        );

    \I__758\ : InMux
    port map (
            O => \N__4616\,
            I => \N__4613\
        );

    \I__757\ : LocalMux
    port map (
            O => \N__4613\,
            I => \N__4610\
        );

    \I__756\ : Span4Mux_h
    port map (
            O => \N__4610\,
            I => \N__4607\
        );

    \I__755\ : Odrv4
    port map (
            O => \N__4607\,
            I => \DFT.multiplier.regsA_un3_result_cry_2_THRU_CO\
        );

    \I__754\ : InMux
    port map (
            O => \N__4604\,
            I => \N__4601\
        );

    \I__753\ : LocalMux
    port map (
            O => \N__4601\,
            I => \N__4598\
        );

    \I__752\ : Span4Mux_v
    port map (
            O => \N__4598\,
            I => \N__4595\
        );

    \I__751\ : Odrv4
    port map (
            O => \N__4595\,
            I => \X_1__10\
        );

    \I__750\ : CascadeMux
    port map (
            O => \N__4592\,
            I => \N__4589\
        );

    \I__749\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4586\
        );

    \I__748\ : LocalMux
    port map (
            O => \N__4586\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_964\
        );

    \I__747\ : InMux
    port map (
            O => \N__4583\,
            I => \DFT.multiplier.regsA_un3_result_cry_2_0\
        );

    \I__746\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4577\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4577\,
            I => \N__4574\
        );

    \I__744\ : Odrv4
    port map (
            O => \N__4574\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_659\
        );

    \I__743\ : InMux
    port map (
            O => \N__4571\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_7\
        );

    \I__742\ : CascadeMux
    port map (
            O => \N__4568\,
            I => \N__4565\
        );

    \I__741\ : InMux
    port map (
            O => \N__4565\,
            I => \N__4562\
        );

    \I__740\ : LocalMux
    port map (
            O => \N__4562\,
            I => \N__4559\
        );

    \I__739\ : Odrv4
    port map (
            O => \N__4559\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_660\
        );

    \I__738\ : InMux
    port map (
            O => \N__4556\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_7\
        );

    \I__737\ : InMux
    port map (
            O => \N__4553\,
            I => \N__4550\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4550\,
            I => \N__4547\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__4547\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_661_THRU_CO\
        );

    \I__734\ : InMux
    port map (
            O => \N__4544\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_661\
        );

    \I__733\ : InMux
    port map (
            O => \N__4541\,
            I => \bfn_11_20_0_\
        );

    \I__732\ : InMux
    port map (
            O => \N__4538\,
            I => \N__4535\
        );

    \I__731\ : LocalMux
    port map (
            O => \N__4535\,
            I => \N__4532\
        );

    \I__730\ : Odrv4
    port map (
            O => \N__4532\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_662_THRU_CO\
        );

    \I__729\ : InMux
    port map (
            O => \N__4529\,
            I => \N__4526\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__4526\,
            I => \N__4523\
        );

    \I__727\ : Odrv4
    port map (
            O => \N__4523\,
            I => \DFT.multiplier.regsA_un3_result_cry_13_0_c_RNO\
        );

    \I__726\ : CascadeMux
    port map (
            O => \N__4520\,
            I => \DFT.state_2_0_cascade_\
        );

    \I__725\ : CascadeMux
    port map (
            O => \N__4517\,
            I => \N__4514\
        );

    \I__724\ : InMux
    port map (
            O => \N__4514\,
            I => \N__4511\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4511\,
            I => \N__4508\
        );

    \I__722\ : Odrv4
    port map (
            O => \N__4508\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_558_THRU_CO\
        );

    \I__721\ : InMux
    port map (
            O => \N__4505\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_558\
        );

    \I__720\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4499\
        );

    \I__719\ : LocalMux
    port map (
            O => \N__4499\,
            I => \N__4496\
        );

    \I__718\ : Odrv4
    port map (
            O => \N__4496\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_559_THRU_CO\
        );

    \I__717\ : InMux
    port map (
            O => \N__4493\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_559\
        );

    \I__716\ : InMux
    port map (
            O => \N__4490\,
            I => \N__4487\
        );

    \I__715\ : LocalMux
    port map (
            O => \N__4487\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_594_THRU_CO\
        );

    \I__714\ : InMux
    port map (
            O => \N__4484\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_560\
        );

    \I__713\ : InMux
    port map (
            O => \N__4481\,
            I => \N__4478\
        );

    \I__712\ : LocalMux
    port map (
            O => \N__4478\,
            I => \N__4475\
        );

    \I__711\ : Odrv4
    port map (
            O => \N__4475\,
            I => \DFT.multiplier.regsA_un3_result_axb_13\
        );

    \I__710\ : CascadeMux
    port map (
            O => \N__4472\,
            I => \N__4469\
        );

    \I__709\ : InMux
    port map (
            O => \N__4469\,
            I => \N__4466\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4466\,
            I => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_3\
        );

    \I__707\ : InMux
    port map (
            O => \N__4463\,
            I => \N__4457\
        );

    \I__706\ : InMux
    port map (
            O => \N__4462\,
            I => \N__4457\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4457\,
            I => \N__4454\
        );

    \I__704\ : Span4Mux_h
    port map (
            O => \N__4454\,
            I => \N__4451\
        );

    \I__703\ : Odrv4
    port map (
            O => \N__4451\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_655_THRU_CO\
        );

    \I__702\ : InMux
    port map (
            O => \N__4448\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_655\
        );

    \I__701\ : InMux
    port map (
            O => \N__4445\,
            I => \N__4442\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4442\,
            I => \N__4439\
        );

    \I__699\ : Odrv4
    port map (
            O => \N__4439\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_656_THRU_CO\
        );

    \I__698\ : InMux
    port map (
            O => \N__4436\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_656\
        );

    \I__697\ : CascadeMux
    port map (
            O => \N__4433\,
            I => \N__4430\
        );

    \I__696\ : InMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__695\ : LocalMux
    port map (
            O => \N__4427\,
            I => \N__4424\
        );

    \I__694\ : Odrv4
    port map (
            O => \N__4424\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_657_THRU_CO\
        );

    \I__693\ : InMux
    port map (
            O => \N__4421\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_657\
        );

    \I__692\ : CascadeMux
    port map (
            O => \N__4418\,
            I => \N__4415\
        );

    \I__691\ : InMux
    port map (
            O => \N__4415\,
            I => \N__4412\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4412\,
            I => \N__4409\
        );

    \I__689\ : Odrv4
    port map (
            O => \N__4409\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_658_THRU_CO\
        );

    \I__688\ : InMux
    port map (
            O => \N__4406\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_658\
        );

    \I__687\ : InMux
    port map (
            O => \N__4403\,
            I => \N__4400\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4400\,
            I => \N__4397\
        );

    \I__685\ : Span4Mux_h
    port map (
            O => \N__4397\,
            I => \N__4394\
        );

    \I__684\ : Odrv4
    port map (
            O => \N__4394\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_550_THRU_CO\
        );

    \I__683\ : InMux
    port map (
            O => \N__4391\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_550\
        );

    \I__682\ : InMux
    port map (
            O => \N__4388\,
            I => \N__4385\
        );

    \I__681\ : LocalMux
    port map (
            O => \N__4385\,
            I => \N__4382\
        );

    \I__680\ : Odrv4
    port map (
            O => \N__4382\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_551\
        );

    \I__679\ : InMux
    port map (
            O => \N__4379\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_6\
        );

    \I__678\ : InMux
    port map (
            O => \N__4376\,
            I => \N__4373\
        );

    \I__677\ : LocalMux
    port map (
            O => \N__4373\,
            I => \N__4370\
        );

    \I__676\ : Span4Mux_h
    port map (
            O => \N__4370\,
            I => \N__4367\
        );

    \I__675\ : Odrv4
    port map (
            O => \N__4367\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_552\
        );

    \I__674\ : InMux
    port map (
            O => \N__4364\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_6\
        );

    \I__673\ : InMux
    port map (
            O => \N__4361\,
            I => \N__4358\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__671\ : Odrv4
    port map (
            O => \N__4355\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_553_THRU_CO\
        );

    \I__670\ : InMux
    port map (
            O => \N__4352\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_553\
        );

    \I__669\ : InMux
    port map (
            O => \N__4349\,
            I => \N__4346\
        );

    \I__668\ : LocalMux
    port map (
            O => \N__4346\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_554_THRU_CO\
        );

    \I__667\ : InMux
    port map (
            O => \N__4343\,
            I => \bfn_11_18_0_\
        );

    \I__666\ : CascadeMux
    port map (
            O => \N__4340\,
            I => \N__4337\
        );

    \I__665\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4334\
        );

    \I__664\ : LocalMux
    port map (
            O => \N__4334\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_555_THRU_CO\
        );

    \I__663\ : InMux
    port map (
            O => \N__4331\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_555\
        );

    \I__662\ : InMux
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4325\,
            I => \N__4322\
        );

    \I__660\ : Span4Mux_h
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__4319\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_556_THRU_CO\
        );

    \I__658\ : InMux
    port map (
            O => \N__4316\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_556\
        );

    \I__657\ : InMux
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__656\ : LocalMux
    port map (
            O => \N__4310\,
            I => \N__4307\
        );

    \I__655\ : Span4Mux_v
    port map (
            O => \N__4307\,
            I => \N__4304\
        );

    \I__654\ : Odrv4
    port map (
            O => \N__4304\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_557_THRU_CO\
        );

    \I__653\ : InMux
    port map (
            O => \N__4301\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_557\
        );

    \I__652\ : InMux
    port map (
            O => \N__4298\,
            I => \N__4295\
        );

    \I__651\ : LocalMux
    port map (
            O => \N__4295\,
            I => \N__4292\
        );

    \I__650\ : Span4Mux_h
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__649\ : Odrv4
    port map (
            O => \N__4289\,
            I => \X_1__11\
        );

    \I__648\ : InMux
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4283\,
            I => \X_1__13\
        );

    \I__646\ : InMux
    port map (
            O => \N__4280\,
            I => \N__4277\
        );

    \I__645\ : LocalMux
    port map (
            O => \N__4277\,
            I => \X_1__12\
        );

    \I__644\ : IoInMux
    port map (
            O => \N__4274\,
            I => \N__4271\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__4271\,
            I => \N__4268\
        );

    \I__642\ : Span12Mux_s8_h
    port map (
            O => \N__4268\,
            I => \N__4265\
        );

    \I__641\ : Odrv12
    port map (
            O => \N__4265\,
            I => \o_X_c_22\
        );

    \I__640\ : IoInMux
    port map (
            O => \N__4262\,
            I => \N__4259\
        );

    \I__639\ : LocalMux
    port map (
            O => \N__4259\,
            I => \N__4256\
        );

    \I__638\ : Span4Mux_s3_h
    port map (
            O => \N__4256\,
            I => \N__4253\
        );

    \I__637\ : Span4Mux_h
    port map (
            O => \N__4253\,
            I => \N__4250\
        );

    \I__636\ : Span4Mux_v
    port map (
            O => \N__4250\,
            I => \N__4247\
        );

    \I__635\ : Odrv4
    port map (
            O => \N__4247\,
            I => \o_X_c_20\
        );

    \I__634\ : InMux
    port map (
            O => \N__4244\,
            I => \N__4241\
        );

    \I__633\ : LocalMux
    port map (
            O => \N__4241\,
            I => \N__4238\
        );

    \I__632\ : Span4Mux_v
    port map (
            O => \N__4238\,
            I => \N__4235\
        );

    \I__631\ : Odrv4
    port map (
            O => \N__4235\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_549_THRU_CO\
        );

    \I__630\ : InMux
    port map (
            O => \N__4232\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_549\
        );

    \I__629\ : InMux
    port map (
            O => \N__4229\,
            I => \N__4226\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__4226\,
            I => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNI8J5C1\
        );

    \I__627\ : CascadeMux
    port map (
            O => \N__4223\,
            I => \N__4219\
        );

    \I__626\ : InMux
    port map (
            O => \N__4222\,
            I => \N__4216\
        );

    \I__625\ : InMux
    port map (
            O => \N__4219\,
            I => \N__4213\
        );

    \I__624\ : LocalMux
    port map (
            O => \N__4216\,
            I => \N__4208\
        );

    \I__623\ : LocalMux
    port map (
            O => \N__4213\,
            I => \N__4208\
        );

    \I__622\ : Odrv4
    port map (
            O => \N__4208\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_825\
        );

    \I__621\ : InMux
    port map (
            O => \N__4205\,
            I => \DFT.multiplier.regsA_un3_result_cry_3_0\
        );

    \I__620\ : InMux
    port map (
            O => \N__4202\,
            I => \N__4199\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4199\,
            I => \N__4196\
        );

    \I__618\ : Odrv4
    port map (
            O => \N__4196\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_826\
        );

    \I__617\ : CascadeMux
    port map (
            O => \N__4193\,
            I => \N__4190\
        );

    \I__616\ : InMux
    port map (
            O => \N__4190\,
            I => \N__4187\
        );

    \I__615\ : LocalMux
    port map (
            O => \N__4187\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_860\
        );

    \I__614\ : InMux
    port map (
            O => \N__4184\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_8\
        );

    \I__613\ : InMux
    port map (
            O => \N__4181\,
            I => \N__4178\
        );

    \I__612\ : LocalMux
    port map (
            O => \N__4178\,
            I => \N__4175\
        );

    \I__611\ : Odrv12
    port map (
            O => \N__4175\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_827\
        );

    \I__610\ : CascadeMux
    port map (
            O => \N__4172\,
            I => \N__4169\
        );

    \I__609\ : InMux
    port map (
            O => \N__4169\,
            I => \N__4166\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__4166\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_861\
        );

    \I__607\ : InMux
    port map (
            O => \N__4163\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_1\
        );

    \I__606\ : InMux
    port map (
            O => \N__4160\,
            I => \N__4157\
        );

    \I__605\ : LocalMux
    port map (
            O => \N__4157\,
            I => \N__4154\
        );

    \I__604\ : Odrv4
    port map (
            O => \N__4154\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_828\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__4151\,
            I => \N__4148\
        );

    \I__602\ : InMux
    port map (
            O => \N__4148\,
            I => \N__4145\
        );

    \I__601\ : LocalMux
    port map (
            O => \N__4145\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_862\
        );

    \I__600\ : InMux
    port map (
            O => \N__4142\,
            I => \DFT.multiplier.regsA_un3_result_cry_6\
        );

    \I__599\ : InMux
    port map (
            O => \N__4139\,
            I => \N__4136\
        );

    \I__598\ : LocalMux
    port map (
            O => \N__4136\,
            I => \N__4133\
        );

    \I__597\ : Odrv12
    port map (
            O => \N__4133\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_829\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__4130\,
            I => \N__4127\
        );

    \I__595\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4124\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__4124\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_863\
        );

    \I__593\ : InMux
    port map (
            O => \N__4121\,
            I => \DFT.multiplier.regsA_un3_result_cry_7\
        );

    \I__592\ : InMux
    port map (
            O => \N__4118\,
            I => \N__4115\
        );

    \I__591\ : LocalMux
    port map (
            O => \N__4115\,
            I => \N__4112\
        );

    \I__590\ : Odrv12
    port map (
            O => \N__4112\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_830\
        );

    \I__589\ : CascadeMux
    port map (
            O => \N__4109\,
            I => \N__4106\
        );

    \I__588\ : InMux
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__587\ : LocalMux
    port map (
            O => \N__4103\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_864\
        );

    \I__586\ : InMux
    port map (
            O => \N__4100\,
            I => \DFT.multiplier.regsA_un3_result_cry_8_0\
        );

    \I__585\ : InMux
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__583\ : Odrv4
    port map (
            O => \N__4091\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_831\
        );

    \I__582\ : CascadeMux
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__581\ : InMux
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__580\ : LocalMux
    port map (
            O => \N__4082\,
            I => \N__4079\
        );

    \I__579\ : Odrv4
    port map (
            O => \N__4079\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_865\
        );

    \I__578\ : InMux
    port map (
            O => \N__4076\,
            I => \bfn_10_23_0_\
        );

    \I__577\ : InMux
    port map (
            O => \N__4073\,
            I => \N__4070\
        );

    \I__576\ : LocalMux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__4067\,
            I => \DFT.multiplier.regsA_un3_result_axb_11\
        );

    \I__574\ : InMux
    port map (
            O => \N__4064\,
            I => \DFT.multiplier.regsA_un3_result_cry_10\
        );

    \I__573\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__571\ : Odrv4
    port map (
            O => \N__4055\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_623\
        );

    \I__570\ : InMux
    port map (
            O => \N__4052\,
            I => \DFT.multiplier.regsA_un3_result_cry_3_2\
        );

    \I__569\ : InMux
    port map (
            O => \N__4049\,
            I => \N__4046\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__567\ : Odrv4
    port map (
            O => \N__4043\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_624\
        );

    \I__566\ : InMux
    port map (
            O => \N__4040\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_1\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__4037\,
            I => \N__4034\
        );

    \I__564\ : InMux
    port map (
            O => \N__4034\,
            I => \N__4031\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4031\,
            I => \N__4028\
        );

    \I__562\ : Odrv4
    port map (
            O => \N__4028\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_625_THRU_CO\
        );

    \I__561\ : InMux
    port map (
            O => \N__4025\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_2\
        );

    \I__560\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4019\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__4019\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_626_THRU_CO\
        );

    \I__558\ : InMux
    port map (
            O => \N__4016\,
            I => \DFT.multiplier.regsA_un3_result_cry_6_0\
        );

    \I__557\ : CascadeMux
    port map (
            O => \N__4013\,
            I => \N__4010\
        );

    \I__556\ : InMux
    port map (
            O => \N__4010\,
            I => \N__4007\
        );

    \I__555\ : LocalMux
    port map (
            O => \N__4007\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_627_THRU_CO\
        );

    \I__554\ : InMux
    port map (
            O => \N__4004\,
            I => \DFT.multiplier.regsA_un3_result_cry_7_0\
        );

    \I__553\ : InMux
    port map (
            O => \N__4001\,
            I => \DFT.multiplier.regsA_un3_result_cry_8\
        );

    \I__552\ : InMux
    port map (
            O => \N__3998\,
            I => \N__3995\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3995\,
            I => \DFT.multiplier.regsA_un3_result_cry_8_THRU_CO\
        );

    \I__550\ : InMux
    port map (
            O => \N__3992\,
            I => \N__3989\
        );

    \I__549\ : LocalMux
    port map (
            O => \N__3989\,
            I => \N__3986\
        );

    \I__548\ : Odrv12
    port map (
            O => \N__3986\,
            I => \X_1__6\
        );

    \I__547\ : InMux
    port map (
            O => \N__3983\,
            I => \N__3980\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3980\,
            I => \N__3977\
        );

    \I__545\ : Span4Mux_h
    port map (
            O => \N__3977\,
            I => \N__3974\
        );

    \I__544\ : Odrv4
    port map (
            O => \N__3974\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_620_THRU_CO\
        );

    \I__543\ : CascadeMux
    port map (
            O => \N__3971\,
            I => \N__3968\
        );

    \I__542\ : InMux
    port map (
            O => \N__3968\,
            I => \N__3965\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3965\,
            I => \N__3962\
        );

    \I__540\ : Odrv12
    port map (
            O => \N__3962\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_824\
        );

    \I__539\ : InMux
    port map (
            O => \N__3959\,
            I => \DFT.multiplier.regsA_un3_result_cry_2_1\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__3956\,
            I => \N__3953\
        );

    \I__537\ : InMux
    port map (
            O => \N__3953\,
            I => \N__3950\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3950\,
            I => \N__3947\
        );

    \I__535\ : Odrv4
    port map (
            O => \N__3947\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_588\
        );

    \I__534\ : InMux
    port map (
            O => \N__3944\,
            I => \DFT.multiplier.regsA_un3_result_cry_6_1\
        );

    \I__533\ : InMux
    port map (
            O => \N__3941\,
            I => \N__3938\
        );

    \I__532\ : LocalMux
    port map (
            O => \N__3938\,
            I => \N__3935\
        );

    \I__531\ : Odrv4
    port map (
            O => \N__3935\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_589_THRU_CO\
        );

    \I__530\ : InMux
    port map (
            O => \N__3932\,
            I => \DFT.multiplier.regsA_un3_result_cry_7_1\
        );

    \I__529\ : CascadeMux
    port map (
            O => \N__3929\,
            I => \N__3926\
        );

    \I__528\ : InMux
    port map (
            O => \N__3926\,
            I => \N__3923\
        );

    \I__527\ : LocalMux
    port map (
            O => \N__3923\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_590_THRU_CO\
        );

    \I__526\ : InMux
    port map (
            O => \N__3920\,
            I => \DFT.multiplier.regsA_un3_result_cry_8_1\
        );

    \I__525\ : CascadeMux
    port map (
            O => \N__3917\,
            I => \N__3914\
        );

    \I__524\ : InMux
    port map (
            O => \N__3914\,
            I => \N__3911\
        );

    \I__523\ : LocalMux
    port map (
            O => \N__3911\,
            I => \N__3908\
        );

    \I__522\ : Odrv4
    port map (
            O => \N__3908\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_591_THRU_CO\
        );

    \I__521\ : InMux
    port map (
            O => \N__3905\,
            I => \bfn_10_20_0_\
        );

    \I__520\ : InMux
    port map (
            O => \N__3902\,
            I => \N__3899\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3899\,
            I => \N__3896\
        );

    \I__518\ : Odrv4
    port map (
            O => \N__3896\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_592_THRU_CO\
        );

    \I__517\ : InMux
    port map (
            O => \N__3893\,
            I => \DFT.multiplier.regsA_un3_result_cry_10_0\
        );

    \I__516\ : CascadeMux
    port map (
            O => \N__3890\,
            I => \N__3887\
        );

    \I__515\ : InMux
    port map (
            O => \N__3887\,
            I => \N__3884\
        );

    \I__514\ : LocalMux
    port map (
            O => \N__3884\,
            I => \N__3881\
        );

    \I__513\ : Odrv4
    port map (
            O => \N__3881\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_593_THRU_CO\
        );

    \I__512\ : InMux
    port map (
            O => \N__3878\,
            I => \DFT.multiplier.regsA_un3_result_cry_11\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__3875\,
            I => \N__3872\
        );

    \I__510\ : InMux
    port map (
            O => \N__3872\,
            I => \N__3869\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3869\,
            I => \DFT.multiplier.regsA_un3_result_axb_9\
        );

    \I__508\ : InMux
    port map (
            O => \N__3866\,
            I => \DFT.multiplier.regsA_un3_result_cry_12\
        );

    \I__507\ : CascadeMux
    port map (
            O => \N__3863\,
            I => \N__3860\
        );

    \I__506\ : InMux
    port map (
            O => \N__3860\,
            I => \N__3857\
        );

    \I__505\ : LocalMux
    port map (
            O => \N__3857\,
            I => \N__3854\
        );

    \I__504\ : Span4Mux_v
    port map (
            O => \N__3854\,
            I => \N__3851\
        );

    \I__503\ : Odrv4
    port map (
            O => \N__3851\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_621_THRU_CO\
        );

    \I__502\ : CascadeMux
    port map (
            O => \N__3848\,
            I => \N__3845\
        );

    \I__501\ : InMux
    port map (
            O => \N__3845\,
            I => \N__3842\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3842\,
            I => \N__3839\
        );

    \I__499\ : Odrv4
    port map (
            O => \N__3839\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_622_THRU_CO\
        );

    \I__498\ : InMux
    port map (
            O => \N__3836\,
            I => \DFT.multiplier.regsA_un3_result_cry_2_3\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__496\ : InMux
    port map (
            O => \N__3830\,
            I => \N__3827\
        );

    \I__495\ : LocalMux
    port map (
            O => \N__3827\,
            I => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_2\
        );

    \I__494\ : CascadeMux
    port map (
            O => \N__3824\,
            I => \N__3821\
        );

    \I__493\ : InMux
    port map (
            O => \N__3821\,
            I => \N__3818\
        );

    \I__492\ : LocalMux
    port map (
            O => \N__3818\,
            I => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_3\
        );

    \I__491\ : CascadeMux
    port map (
            O => \N__3815\,
            I => \N__3812\
        );

    \I__490\ : InMux
    port map (
            O => \N__3812\,
            I => \N__3809\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3809\,
            I => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_2\
        );

    \I__488\ : CascadeMux
    port map (
            O => \N__3806\,
            I => \N__3803\
        );

    \I__487\ : InMux
    port map (
            O => \N__3803\,
            I => \N__3800\
        );

    \I__486\ : LocalMux
    port map (
            O => \N__3800\,
            I => \N__3797\
        );

    \I__485\ : Odrv4
    port map (
            O => \N__3797\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_583_THRU_CO\
        );

    \I__484\ : CascadeMux
    port map (
            O => \N__3794\,
            I => \N__3791\
        );

    \I__483\ : InMux
    port map (
            O => \N__3791\,
            I => \N__3788\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3788\,
            I => \N__3785\
        );

    \I__481\ : Odrv4
    port map (
            O => \N__3785\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_584_THRU_CO\
        );

    \I__480\ : CascadeMux
    port map (
            O => \N__3782\,
            I => \N__3779\
        );

    \I__479\ : InMux
    port map (
            O => \N__3779\,
            I => \N__3776\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3776\,
            I => \N__3773\
        );

    \I__477\ : Odrv4
    port map (
            O => \N__3773\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_585_THRU_CO\
        );

    \I__476\ : InMux
    port map (
            O => \N__3770\,
            I => \DFT.multiplier.regsA_un3_result_cry_3_3\
        );

    \I__475\ : CascadeMux
    port map (
            O => \N__3767\,
            I => \N__3764\
        );

    \I__474\ : InMux
    port map (
            O => \N__3764\,
            I => \N__3761\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3761\,
            I => \N__3758\
        );

    \I__472\ : Odrv12
    port map (
            O => \N__3758\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_586_THRU_CO\
        );

    \I__471\ : InMux
    port map (
            O => \N__3755\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_2\
        );

    \I__470\ : CascadeMux
    port map (
            O => \N__3752\,
            I => \N__3749\
        );

    \I__469\ : InMux
    port map (
            O => \N__3749\,
            I => \N__3746\
        );

    \I__468\ : LocalMux
    port map (
            O => \N__3746\,
            I => \N__3743\
        );

    \I__467\ : Odrv4
    port map (
            O => \N__3743\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_587\
        );

    \I__466\ : InMux
    port map (
            O => \N__3740\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_3\
        );

    \I__465\ : InMux
    port map (
            O => \N__3737\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_586\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__3734\,
            I => \N__3731\
        );

    \I__463\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3728\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_ma_1\
        );

    \I__461\ : InMux
    port map (
            O => \N__3725\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_5\
        );

    \I__460\ : InMux
    port map (
            O => \N__3722\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_5\
        );

    \I__459\ : InMux
    port map (
            O => \N__3719\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_589\
        );

    \I__458\ : InMux
    port map (
            O => \N__3716\,
            I => \bfn_10_18_0_\
        );

    \I__457\ : InMux
    port map (
            O => \N__3713\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_591\
        );

    \I__456\ : InMux
    port map (
            O => \N__3710\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_592\
        );

    \I__455\ : InMux
    port map (
            O => \N__3707\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_593\
        );

    \I__454\ : InMux
    port map (
            O => \N__3704\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_594\
        );

    \I__453\ : InMux
    port map (
            O => \N__3701\,
            I => \N__3698\
        );

    \I__452\ : LocalMux
    port map (
            O => \N__3698\,
            I => \N__3695\
        );

    \I__451\ : Odrv4
    port map (
            O => \N__3695\,
            I => \X_1__8\
        );

    \I__450\ : InMux
    port map (
            O => \N__3692\,
            I => \N__3689\
        );

    \I__449\ : LocalMux
    port map (
            O => \N__3689\,
            I => \N__3686\
        );

    \I__448\ : Odrv4
    port map (
            O => \N__3686\,
            I => \X_1__9\
        );

    \I__447\ : InMux
    port map (
            O => \N__3683\,
            I => \N__3680\
        );

    \I__446\ : LocalMux
    port map (
            O => \N__3680\,
            I => \X_1__7\
        );

    \I__445\ : IoInMux
    port map (
            O => \N__3677\,
            I => \N__3674\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3674\,
            I => \N__3671\
        );

    \I__443\ : Span4Mux_s0_v
    port map (
            O => \N__3671\,
            I => \N__3668\
        );

    \I__442\ : Sp12to4
    port map (
            O => \N__3668\,
            I => \N__3665\
        );

    \I__441\ : Span12Mux_s8_h
    port map (
            O => \N__3665\,
            I => \N__3662\
        );

    \I__440\ : Odrv12
    port map (
            O => \N__3662\,
            I => \o_X_c_17\
        );

    \I__439\ : IoInMux
    port map (
            O => \N__3659\,
            I => \N__3656\
        );

    \I__438\ : LocalMux
    port map (
            O => \N__3656\,
            I => \N__3653\
        );

    \I__437\ : IoSpan4Mux
    port map (
            O => \N__3653\,
            I => \N__3650\
        );

    \I__436\ : Span4Mux_s3_h
    port map (
            O => \N__3650\,
            I => \N__3647\
        );

    \I__435\ : Span4Mux_h
    port map (
            O => \N__3647\,
            I => \N__3644\
        );

    \I__434\ : Odrv4
    port map (
            O => \N__3644\,
            I => \o_X_c_23\
        );

    \I__433\ : InMux
    port map (
            O => \N__3641\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_583\
        );

    \I__432\ : InMux
    port map (
            O => \N__3638\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_584\
        );

    \I__431\ : InMux
    port map (
            O => \N__3635\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_585\
        );

    \I__430\ : CascadeMux
    port map (
            O => \N__3632\,
            I => \N__3629\
        );

    \I__429\ : InMux
    port map (
            O => \N__3629\,
            I => \N__3626\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3626\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_0\
        );

    \I__427\ : InMux
    port map (
            O => \N__3623\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_622\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__3620\,
            I => \N__3617\
        );

    \I__425\ : InMux
    port map (
            O => \N__3617\,
            I => \N__3614\
        );

    \I__424\ : LocalMux
    port map (
            O => \N__3614\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_ma_0\
        );

    \I__423\ : InMux
    port map (
            O => \N__3611\,
            I => \DFT.multiplier.regsA_un3_result_cry_4_4\
        );

    \I__422\ : InMux
    port map (
            O => \N__3608\,
            I => \DFT.multiplier.regsA_un3_result_cry_5_4\
        );

    \I__421\ : InMux
    port map (
            O => \N__3605\,
            I => \N__3602\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3602\,
            I => \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO\
        );

    \I__419\ : InMux
    port map (
            O => \N__3599\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_625\
        );

    \I__418\ : InMux
    port map (
            O => \N__3596\,
            I => \bfn_9_20_0_\
        );

    \I__417\ : InMux
    port map (
            O => \N__3593\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_627\
        );

    \I__416\ : InMux
    port map (
            O => \N__3590\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_628\
        );

    \I__415\ : InMux
    port map (
            O => \N__3587\,
            I => \N__3584\
        );

    \I__414\ : LocalMux
    port map (
            O => \N__3584\,
            I => \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO\
        );

    \I__413\ : InMux
    port map (
            O => \N__3581\,
            I => \N__3578\
        );

    \I__412\ : LocalMux
    port map (
            O => \N__3578\,
            I => \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO\
        );

    \I__411\ : CascadeMux
    port map (
            O => \N__3575\,
            I => \N__3572\
        );

    \I__410\ : InMux
    port map (
            O => \N__3572\,
            I => \N__3569\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3569\,
            I => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_2\
        );

    \I__408\ : CascadeMux
    port map (
            O => \N__3566\,
            I => \N__3563\
        );

    \I__407\ : InMux
    port map (
            O => \N__3563\,
            I => \N__3560\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3560\,
            I => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_2\
        );

    \I__405\ : InMux
    port map (
            O => \N__3557\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_619\
        );

    \I__404\ : CascadeMux
    port map (
            O => \N__3554\,
            I => \N__3551\
        );

    \I__403\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3548\
        );

    \I__402\ : LocalMux
    port map (
            O => \N__3548\,
            I => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_1\
        );

    \I__401\ : InMux
    port map (
            O => \N__3545\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_620\
        );

    \I__400\ : CascadeMux
    port map (
            O => \N__3542\,
            I => \N__3539\
        );

    \I__399\ : InMux
    port map (
            O => \N__3539\,
            I => \N__3536\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3536\,
            I => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_1\
        );

    \I__397\ : InMux
    port map (
            O => \N__3533\,
            I => \DFT.multiplier.mult1_AdderTree2i_bigtree_621\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__3530\,
            I => \DFT.o_done_RNOZ0Z_0_cascade_\
        );

    \I__395\ : IoInMux
    port map (
            O => \N__3527\,
            I => \N__3524\
        );

    \I__394\ : LocalMux
    port map (
            O => \N__3524\,
            I => \N__3521\
        );

    \I__393\ : IoSpan4Mux
    port map (
            O => \N__3521\,
            I => \N__3518\
        );

    \I__392\ : IoSpan4Mux
    port map (
            O => \N__3518\,
            I => \N__3515\
        );

    \I__391\ : IoSpan4Mux
    port map (
            O => \N__3515\,
            I => \N__3511\
        );

    \I__390\ : InMux
    port map (
            O => \N__3514\,
            I => \N__3508\
        );

    \I__389\ : IoSpan4Mux
    port map (
            O => \N__3511\,
            I => \N__3505\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3508\,
            I => \N__3502\
        );

    \I__387\ : Span4Mux_s1_h
    port map (
            O => \N__3505\,
            I => \N__3496\
        );

    \I__386\ : Span4Mux_v
    port map (
            O => \N__3502\,
            I => \N__3496\
        );

    \I__385\ : InMux
    port map (
            O => \N__3501\,
            I => \N__3493\
        );

    \I__384\ : Span4Mux_h
    port map (
            O => \N__3496\,
            I => \N__3490\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3493\,
            I => done_c
        );

    \I__382\ : Odrv4
    port map (
            O => \N__3490\,
            I => done_c
        );

    \I__381\ : InMux
    port map (
            O => \N__3485\,
            I => \N__3482\
        );

    \I__380\ : LocalMux
    port map (
            O => \N__3482\,
            I => \N__3478\
        );

    \I__379\ : InMux
    port map (
            O => \N__3481\,
            I => \N__3475\
        );

    \I__378\ : Odrv4
    port map (
            O => \N__3478\,
            I => \DFT.state_RNIHM3GZ0Z_0\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3475\,
            I => \DFT.state_RNIHM3GZ0Z_0\
        );

    \I__376\ : IoInMux
    port map (
            O => \N__3470\,
            I => \N__3467\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__3467\,
            I => \N__3464\
        );

    \I__374\ : IoSpan4Mux
    port map (
            O => \N__3464\,
            I => \N__3461\
        );

    \I__373\ : Span4Mux_s2_h
    port map (
            O => \N__3461\,
            I => \N__3458\
        );

    \I__372\ : Span4Mux_h
    port map (
            O => \N__3458\,
            I => \N__3455\
        );

    \I__371\ : Odrv4
    port map (
            O => \N__3455\,
            I => \o_X_c_18\
        );

    \I__370\ : IoInMux
    port map (
            O => \N__3452\,
            I => \N__3449\
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3449\,
            I => \N__3446\
        );

    \I__368\ : IoSpan4Mux
    port map (
            O => \N__3446\,
            I => \N__3443\
        );

    \I__367\ : Span4Mux_s3_v
    port map (
            O => \N__3443\,
            I => \N__3440\
        );

    \I__366\ : Span4Mux_v
    port map (
            O => \N__3440\,
            I => \N__3437\
        );

    \I__365\ : Odrv4
    port map (
            O => \N__3437\,
            I => \o_X_c_16\
        );

    \I__364\ : IoInMux
    port map (
            O => \N__3434\,
            I => \N__3431\
        );

    \I__363\ : LocalMux
    port map (
            O => \N__3431\,
            I => \N__3428\
        );

    \I__362\ : Span4Mux_s3_h
    port map (
            O => \N__3428\,
            I => \N__3425\
        );

    \I__361\ : Span4Mux_v
    port map (
            O => \N__3425\,
            I => \N__3422\
        );

    \I__360\ : Odrv4
    port map (
            O => \N__3422\,
            I => \o_X_c_19\
        );

    \I__359\ : IoInMux
    port map (
            O => \N__3419\,
            I => \N__3416\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3416\,
            I => \N__3413\
        );

    \I__357\ : IoSpan4Mux
    port map (
            O => \N__3413\,
            I => \N__3410\
        );

    \I__356\ : Span4Mux_s2_h
    port map (
            O => \N__3410\,
            I => \N__3407\
        );

    \I__355\ : Span4Mux_h
    port map (
            O => \N__3407\,
            I => \N__3404\
        );

    \I__354\ : Odrv4
    port map (
            O => \N__3404\,
            I => \o_X_c_21\
        );

    \I__353\ : IoInMux
    port map (
            O => \N__3401\,
            I => \N__3398\
        );

    \I__352\ : LocalMux
    port map (
            O => \N__3398\,
            I => \N__3395\
        );

    \I__351\ : IoSpan4Mux
    port map (
            O => \N__3395\,
            I => \N__3392\
        );

    \I__350\ : Span4Mux_s1_v
    port map (
            O => \N__3392\,
            I => \N__3389\
        );

    \I__349\ : Sp12to4
    port map (
            O => \N__3389\,
            I => \N__3386\
        );

    \I__348\ : Span12Mux_s9_v
    port map (
            O => \N__3386\,
            I => \N__3383\
        );

    \I__347\ : Span12Mux_v
    port map (
            O => \N__3383\,
            I => \N__3380\
        );

    \I__346\ : Odrv12
    port map (
            O => \N__3380\,
            I => i_ref_clk_c
        );

    \I__345\ : IoInMux
    port map (
            O => \N__3377\,
            I => \N__3374\
        );

    \I__344\ : LocalMux
    port map (
            O => \N__3374\,
            I => i_rst_c_i
        );

    \I__343\ : IoInMux
    port map (
            O => \N__3371\,
            I => \N__3368\
        );

    \I__342\ : LocalMux
    port map (
            O => \N__3368\,
            I => \DFT.done_c_0\
        );

    \I__341\ : ClkMux
    port map (
            O => \N__3365\,
            I => \N__3278\
        );

    \I__340\ : ClkMux
    port map (
            O => \N__3364\,
            I => \N__3278\
        );

    \I__339\ : ClkMux
    port map (
            O => \N__3363\,
            I => \N__3278\
        );

    \I__338\ : ClkMux
    port map (
            O => \N__3362\,
            I => \N__3278\
        );

    \I__337\ : ClkMux
    port map (
            O => \N__3361\,
            I => \N__3278\
        );

    \I__336\ : ClkMux
    port map (
            O => \N__3360\,
            I => \N__3278\
        );

    \I__335\ : ClkMux
    port map (
            O => \N__3359\,
            I => \N__3278\
        );

    \I__334\ : ClkMux
    port map (
            O => \N__3358\,
            I => \N__3278\
        );

    \I__333\ : ClkMux
    port map (
            O => \N__3357\,
            I => \N__3278\
        );

    \I__332\ : ClkMux
    port map (
            O => \N__3356\,
            I => \N__3278\
        );

    \I__331\ : ClkMux
    port map (
            O => \N__3355\,
            I => \N__3278\
        );

    \I__330\ : ClkMux
    port map (
            O => \N__3354\,
            I => \N__3278\
        );

    \I__329\ : ClkMux
    port map (
            O => \N__3353\,
            I => \N__3278\
        );

    \I__328\ : ClkMux
    port map (
            O => \N__3352\,
            I => \N__3278\
        );

    \I__327\ : ClkMux
    port map (
            O => \N__3351\,
            I => \N__3278\
        );

    \I__326\ : ClkMux
    port map (
            O => \N__3350\,
            I => \N__3278\
        );

    \I__325\ : ClkMux
    port map (
            O => \N__3349\,
            I => \N__3278\
        );

    \I__324\ : ClkMux
    port map (
            O => \N__3348\,
            I => \N__3278\
        );

    \I__323\ : ClkMux
    port map (
            O => \N__3347\,
            I => \N__3278\
        );

    \I__322\ : ClkMux
    port map (
            O => \N__3346\,
            I => \N__3278\
        );

    \I__321\ : ClkMux
    port map (
            O => \N__3345\,
            I => \N__3278\
        );

    \I__320\ : ClkMux
    port map (
            O => \N__3344\,
            I => \N__3278\
        );

    \I__319\ : ClkMux
    port map (
            O => \N__3343\,
            I => \N__3278\
        );

    \I__318\ : ClkMux
    port map (
            O => \N__3342\,
            I => \N__3278\
        );

    \I__317\ : ClkMux
    port map (
            O => \N__3341\,
            I => \N__3278\
        );

    \I__316\ : ClkMux
    port map (
            O => \N__3340\,
            I => \N__3278\
        );

    \I__315\ : ClkMux
    port map (
            O => \N__3339\,
            I => \N__3278\
        );

    \I__314\ : ClkMux
    port map (
            O => \N__3338\,
            I => \N__3278\
        );

    \I__313\ : ClkMux
    port map (
            O => \N__3337\,
            I => \N__3278\
        );

    \I__312\ : GlobalMux
    port map (
            O => \N__3278\,
            I => \N__3275\
        );

    \I__311\ : gio2CtrlBuf
    port map (
            O => \N__3275\,
            I => sys_clk_g
        );

    \I__310\ : IoInMux
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__309\ : LocalMux
    port map (
            O => \N__3269\,
            I => \N__3266\
        );

    \I__308\ : Odrv4
    port map (
            O => \N__3266\,
            I => sys_clk
        );

    \INVo_X_0__nesr_5C\ : INV
    port map (
            O => \INVo_X_0__nesr_5C_net\,
            I => \N__3338\
        );

    \INVo_X_1__nesr_9C\ : INV
    port map (
            O => \INVo_X_1__nesr_9C_net\,
            I => \N__3342\
        );

    \INVo_X_0__nesr_8C\ : INV
    port map (
            O => \INVo_X_0__nesr_8C_net\,
            I => \N__3339\
        );

    \INVo_X_0__nesr_4C\ : INV
    port map (
            O => \INVo_X_0__nesr_4C_net\,
            I => \N__3341\
        );

    \INVo_X_0__nesr_3C\ : INV
    port map (
            O => \INVo_X_0__nesr_3C_net\,
            I => \N__3348\
        );

    \INVo_X_1__nesr_8C\ : INV
    port map (
            O => \INVo_X_1__nesr_8C_net\,
            I => \N__3352\
        );

    \INVo_X_0__nesr_1C\ : INV
    port map (
            O => \INVo_X_0__nesr_1C_net\,
            I => \N__3354\
        );

    \INVo_X_0__nesr_7C\ : INV
    port map (
            O => \INVo_X_0__nesr_7C_net\,
            I => \N__3337\
        );

    \INVDFT.o_X_0__nesr_6C\ : INV
    port map (
            O => \INVDFT.o_X_0__nesr_6C_net\,
            I => \N__3353\
        );

    \INVDFT.o_X_0__nesr_11C\ : INV
    port map (
            O => \INVDFT.o_X_0__nesr_11C_net\,
            I => \N__3344\
        );

    \INVDFT.o_X_0__nesr_14C\ : INV
    port map (
            O => \INVDFT.o_X_0__nesr_14C_net\,
            I => \N__3347\
        );

    \INVDFT.o_X_0__nesr_10C\ : INV
    port map (
            O => \INVDFT.o_X_0__nesr_10C_net\,
            I => \N__3351\
        );

    \INVDFT.b_6C\ : INV
    port map (
            O => \INVDFT.b_6C_net\,
            I => \N__3362\
        );

    \INVo_X_0__nesr_9C\ : INV
    port map (
            O => \INVo_X_0__nesr_9C_net\,
            I => \N__3340\
        );

    \INVDFT.o_X_0__nesr_13C\ : INV
    port map (
            O => \INVDFT.o_X_0__nesr_13C_net\,
            I => \N__3346\
        );

    \INVDFT.o_X_1__nesr_10C\ : INV
    port map (
            O => \INVDFT.o_X_1__nesr_10C_net\,
            I => \N__3350\
        );

    \INVDFT.o_X_0__nesr_7C\ : INV
    port map (
            O => \INVDFT.o_X_0__nesr_7C_net\,
            I => \N__3357\
        );

    \INVDFT.state_0C\ : INV
    port map (
            O => \INVDFT.state_0C_net\,
            I => \N__3360\
        );

    \INVo_X_1__nesr_4C\ : INV
    port map (
            O => \INVo_X_1__nesr_4C_net\,
            I => \N__3343\
        );

    \INVo_X_1__nesr_6C\ : INV
    port map (
            O => \INVo_X_1__nesr_6C_net\,
            I => \N__3345\
        );

    \INVDFT.o_X_1__nesr_12C\ : INV
    port map (
            O => \INVDFT.o_X_1__nesr_12C_net\,
            I => \N__3349\
        );

    \INVDFT.o_X_1__nesr_6C\ : INV
    port map (
            O => \INVDFT.o_X_1__nesr_6C_net\,
            I => \N__3356\
        );

    \INVo_X_1__nesr_1C\ : INV
    port map (
            O => \INVo_X_1__nesr_1C_net\,
            I => \N__3355\
        );

    \INVDFT.o_X_1__nesr_7C\ : INV
    port map (
            O => \INVDFT.o_X_1__nesr_7C_net\,
            I => \N__3359\
        );

    \INVDFT.o_X_1__nesr_8C\ : INV
    port map (
            O => \INVDFT.o_X_1__nesr_8C_net\,
            I => \N__3361\
        );

    \INVo_X_1__nesr_5C\ : INV
    port map (
            O => \INVo_X_1__nesr_5C_net\,
            I => \N__3358\
        );

    \INVo_X_1__nesr_3C\ : INV
    port map (
            O => \INVo_X_1__nesr_3C_net\,
            I => \N__3363\
        );

    \INVo_X_1__nesr_2C\ : INV
    port map (
            O => \INVo_X_1__nesr_2C_net\,
            I => \N__3364\
        );

    \INVDFT.o_doneC\ : INV
    port map (
            O => \INVDFT.o_doneC_net\,
            I => \N__3365\
        );

    \IN_MUX_bfv_10_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_19_0_\
        );

    \IN_MUX_bfv_10_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DFT.multiplier.regsA_un3_result_cry_9_0\,
            carryinitout => \bfn_10_20_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_14_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_17_0_\
        );

    \IN_MUX_bfv_14_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_14_18_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_11_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DFT.multiplier.mult1_AdderTree2i_bigtree_662\,
            carryinitout => \bfn_11_20_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_9_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DFT.multiplier.mult1_AdderTree2i_bigtree_626\,
            carryinitout => \bfn_9_20_0_\
        );

    \IN_MUX_bfv_10_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_17_0_\
        );

    \IN_MUX_bfv_10_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DFT.multiplier.mult1_AdderTree2i_bigtree_590\,
            carryinitout => \bfn_10_18_0_\
        );

    \IN_MUX_bfv_11_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_17_0_\
        );

    \IN_MUX_bfv_11_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DFT.multiplier.mult1_AdderTree2i_bigtree_554\,
            carryinitout => \bfn_11_18_0_\
        );

    \IN_MUX_bfv_11_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_22_0_\
        );

    \IN_MUX_bfv_13_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_17_0_\
        );

    \IN_MUX_bfv_11_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_23_0_\
        );

    \IN_MUX_bfv_10_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_21_0_\
        );

    \IN_MUX_bfv_10_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_10_22_0_\
        );

    \IN_MUX_bfv_10_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DFT.multiplier.regsA_un3_result_cry_9\,
            carryinitout => \bfn_10_23_0_\
        );

    \DFT.o_done_RNI6TUH_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3371\,
            GLOBALBUFFEROUTPUT => done_c_0_g
        );

    \sys_clk_derived_clock_RNI5LTF\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3272\,
            GLOBALBUFFEROUTPUT => sys_clk_g
        );

    \i_rst_ibuf_RNI6EKC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3377\,
            GLOBALBUFFEROUTPUT => i_rst_c_i_g
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \i_rst_ibuf_RNI6EKC_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__5186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => i_rst_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.o_done_RNI6TUH_LC_1_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__6528\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3514\,
            lcout => \DFT.done_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.o_done_RNO_0_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110111"
        )
    port map (
            in0 => \N__5179\,
            in1 => \N__5222\,
            in2 => \_gnd_net_\,
            in3 => \N__5078\,
            lcout => OPEN,
            ltout => \DFT.o_done_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.o_done_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3485\,
            in2 => \N__3530\,
            in3 => \N__3501\,
            lcout => done_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_doneC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.state_RNIHM3G_0_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__5178\,
            in1 => \N__5217\,
            in2 => \_gnd_net_\,
            in3 => \N__5072\,
            lcout => \DFT.state_RNIHM3GZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.state_RNIN4OS_0_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6529\,
            in2 => \_gnd_net_\,
            in3 => \N__3481\,
            lcout => \DFT.un1_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_X_1__nesr_2_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3701\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \o_X_c_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_1__nesr_2C_net\,
            ce => \N__6567\,
            sr => \N__6490\
        );

    \o_X_1__nesr_0_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3992\,
            lcout => \o_X_c_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_1__nesr_2C_net\,
            ce => \N__6567\,
            sr => \N__6490\
        );

    \o_X_1__nesr_3_LC_7_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3692\,
            lcout => \o_X_c_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_1__nesr_3C_net\,
            ce => \N__6568\,
            sr => \N__6491\
        );

    \o_X_1__nesr_5_LC_7_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4298\,
            lcout => \o_X_c_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_1__nesr_5C_net\,
            ce => \N__6569\,
            sr => \N__6498\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_1_0_c_RNO_LC_9_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5929\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_4_0_c_RNO_LC_9_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5933\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_7_0_c_RNO_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5935\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_5_ma_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5934\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_5_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_2_0_c_RNO_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5931\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_5_ma_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5930\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_5_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_3_0_c_RNO_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5932\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_0_0_c_RNO_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5928\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_0_0_c_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3575\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_619\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_LUT4_0_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3566\,
            in3 => \N__3557\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_619\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_620\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_620_THRU_LUT4_0_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3554\,
            in3 => \N__3545\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_620_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_620\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_621\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_621_THRU_LUT4_0_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3542\,
            in3 => \N__3533\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_621_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_621\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_622\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_622_THRU_LUT4_0_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3632\,
            in3 => \N__3623\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_622_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_622\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_4_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_4_0_c_RNIHHTP_LC_9_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6044\,
            in2 => \N__3620\,
            in3 => \N__3611\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_623\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_4_4\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_5_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_5_0_c_RNITTRA_LC_9_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5969\,
            in3 => \N__3608\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_624\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_5_4\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_625\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_625_THRU_LUT4_0_LC_9_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3605\,
            in2 => \_gnd_net_\,
            in3 => \N__3599\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_625_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_625\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_626\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_626_THRU_LUT4_0_LC_9_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3587\,
            in2 => \_gnd_net_\,
            in3 => \N__3596\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_626_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_9_20_0_\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_627\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_627_THRU_LUT4_0_LC_9_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3581\,
            in2 => \_gnd_net_\,
            in3 => \N__3593\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_627_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_627\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_628\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_7_0_c_RNIVTM7_LC_9_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4538\,
            in2 => \_gnd_net_\,
            in3 => \N__3590\,
            lcout => \DFT.multiplier.regsA_un3_result_axb_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_8_0_c_RNO_LC_9_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5952\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_9_0_c_RNO_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5953\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.o_X_1__nesr_8_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4633\,
            lcout => \X_1__8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_1__nesr_8C_net\,
            ce => \N__4750\,
            sr => \N__6495\
        );

    \DFT.o_X_1__nesr_7_LC_9_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4658\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \X_1__7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_1__nesr_7C_net\,
            ce => \N__4758\,
            sr => \N__6499\
        );

    \DFT.o_X_1__nesr_9_LC_9_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4646\,
            lcout => \X_1__9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_1__nesr_7C_net\,
            ce => \N__4758\,
            sr => \N__6499\
        );

    \o_X_1__nesr_1_LC_9_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3683\,
            lcout => \o_X_c_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_1__nesr_1C_net\,
            ce => \N__6571\,
            sr => \N__6502\
        );

    \o_X_1__nesr_7_LC_9_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4286\,
            lcout => \o_X_c_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_1__nesr_1C_net\,
            ce => \N__6571\,
            sr => \N__6502\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_0_0_c_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4472\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_17_0_\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_583\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_583_THRU_LUT4_0_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3824\,
            in3 => \N__3641\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_583_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_583\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_584\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_584_THRU_LUT4_0_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3815\,
            in3 => \N__3638\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_584_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_584\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_585\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_585_THRU_LUT4_0_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3833\,
            in3 => \N__3635\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_585_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_585\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_586\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_586_THRU_LUT4_0_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4856\,
            in3 => \N__3737\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_586_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_586\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_4_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_4_0_c_RNIGMTH_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5402\,
            in2 => \N__3734\,
            in3 => \N__3725\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_587\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_4_5\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_5_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_5_0_c_RNIS2SI_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5393\,
            in3 => \N__3722\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_588\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_5_5\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_589\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_589_THRU_LUT4_0_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5414\,
            in3 => \N__3719\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_589_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_589\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_590\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_590_THRU_LUT4_0_LC_10_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5702\,
            in3 => \N__3716\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_590_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_10_18_0_\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_591\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_591_THRU_LUT4_0_LC_10_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5510\,
            in2 => \_gnd_net_\,
            in3 => \N__3713\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_591_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_591\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_592\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_592_THRU_LUT4_0_LC_10_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5000\,
            in2 => \_gnd_net_\,
            in3 => \N__3710\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_592_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_592\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_593\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_593_THRU_LUT4_0_LC_10_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4670\,
            in2 => \_gnd_net_\,
            in3 => \N__3707\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_593_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_593\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_594\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_594_THRU_LUT4_0_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3704\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_594_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_3_0_c_RNO_LC_10_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5927\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_1_0_c_RNO_LC_10_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5925\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_2_0_c_RNO_LC_10_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5926\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_2_c_LC_10_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4244\,
            in2 => \N__3806\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_10_19_0_\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_2_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_3_c_LC_10_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4403\,
            in2 => \N__3794\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_2_4\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_3_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIS12B1_LC_10_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4388\,
            in2 => \N__3782\,
            in3 => \N__3770\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_823\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_3_3\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_4_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNIK3NM_LC_10_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4376\,
            in2 => \N__3767\,
            in3 => \N__3755\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_824\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_4_2\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_5_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIND4V_LC_10_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4361\,
            in2 => \N__3752\,
            in3 => \N__3740\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_825\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_5_3\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_6_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNI50A41_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4349\,
            in2 => \N__3956\,
            in3 => \N__3944\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_826\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_6_1\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_7_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_7_c_RNINH451_LC_10_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3941\,
            in2 => \N__4340\,
            in3 => \N__3932\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_827\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_7_1\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_8_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_8_c_RNIQRHD_LC_10_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4328\,
            in2 => \N__3929\,
            in3 => \N__3920\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_828\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_8_1\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_9_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_9_c_RNI4O6E_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4313\,
            in2 => \N__3917\,
            in3 => \N__3905\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_829\,
            ltout => OPEN,
            carryin => \bfn_10_20_0_\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_10_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_10_c_RNIE7KN_LC_10_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3902\,
            in2 => \N__4517\,
            in3 => \N__3893\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_830\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_10_0\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_11_c_RNIO44O_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4502\,
            in2 => \N__3890\,
            in3 => \N__3878\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_831\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_11\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_12_c_RNIQFFJ1_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__4481\,
            in1 => \N__3998\,
            in2 => \N__3875\,
            in3 => \N__3866\,
            lcout => \DFT.multiplier.regsA_un3_result_axb_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_RNI8J5C1_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__4222\,
            in1 => \N__4462\,
            in2 => \N__3863\,
            in3 => \N__4463\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNI8J5C1\,
            ltout => OPEN,
            carryin => \bfn_10_21_0_\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_2_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_2_c_RNID4E01_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4445\,
            in2 => \N__3848\,
            in3 => \N__3836\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_860\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_2_3\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_3_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_3_c_RNIMULJ1_LC_10_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4061\,
            in2 => \N__4433\,
            in3 => \N__4052\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_861\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_3_2\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_4_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_4_c_RNI4HRO_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4049\,
            in2 => \N__4418\,
            in3 => \N__4040\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_862\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_4_1\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_5_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_5_c_RNISIG41_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4580\,
            in2 => \N__4037\,
            in3 => \N__4025\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_863\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_5_2\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_6_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_6_c_RNIA5M91_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4022\,
            in2 => \N__4568\,
            in3 => \N__4016\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_864\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_6_0\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_7_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_7_c_RNISMGA1_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4553\,
            in2 => \N__4013\,
            in3 => \N__4004\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_865\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_7_0\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.regsA_un3_result_cry_8_THRU_LUT4_0_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4001\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.o_X_1__nesr_6_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5686\,
            in2 => \N__5662\,
            in3 => \_gnd_net_\,
            lcout => \X_1__6\,
            ltout => OPEN,
            carryin => \bfn_10_22_0_\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_2_1\,
            clk => \INVDFT.o_X_1__nesr_6C_net\,
            ce => \N__4751\,
            sr => \N__6496\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_2_c_RNIMU8V_LC_10_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3983\,
            in2 => \N__3971\,
            in3 => \N__3959\,
            lcout => \DFT.x_7\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_2_1\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_3_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIQ8CH2_LC_10_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4229\,
            in2 => \N__4223\,
            in3 => \N__4205\,
            lcout => \DFT.x_8\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_3_0\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_4_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNIEERA2_LC_10_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4202\,
            in2 => \N__4193\,
            in3 => \N__4184\,
            lcout => \DFT.x_9\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_4_8\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_5_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIASUU2_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4181\,
            in2 => \N__4172\,
            in3 => \N__4163\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_963\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_5_1\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNISQIC1_LC_10_22_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4160\,
            in2 => \N__4151\,
            in3 => \N__4142\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_964\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_6\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_7_c_RNIVQTO1_LC_10_22_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4139\,
            in2 => \N__4130\,
            in3 => \N__4121\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_965\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_7\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_8_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_8_c_RNIOUH72_LC_10_22_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4118\,
            in2 => \N__4109\,
            in3 => \N__4100\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_966\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_8_0\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_9_c_RNILFT82_LC_10_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4097\,
            in2 => \N__4088\,
            in3 => \N__4076\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_967\,
            ltout => OPEN,
            carryin => \bfn_10_23_0_\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_10_c_RNITHMQ2_LC_10_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__5378\,
            in1 => \N__4073\,
            in2 => \N__4619\,
            in3 => \N__4064\,
            lcout => \DFT.multiplier.regsA_un3_result_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.o_X_1__nesr_12_LC_10_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4694\,
            lcout => \X_1__12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_1__nesr_12C_net\,
            ce => \N__4763\,
            sr => \N__6503\
        );

    \DFT.o_X_1__nesr_11_LC_10_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5312\,
            in3 => \_gnd_net_\,
            lcout => \X_1__11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_1__nesr_12C_net\,
            ce => \N__4763\,
            sr => \N__6503\
        );

    \DFT.o_X_1__nesr_13_LC_10_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4706\,
            lcout => \X_1__13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_1__nesr_12C_net\,
            ce => \N__4763\,
            sr => \N__6503\
        );

    \o_X_1__nesr_6_LC_10_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4280\,
            lcout => \o_X_c_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_1__nesr_6C_net\,
            ce => \N__6573\,
            sr => \N__6507\
        );

    \o_X_1__nesr_4_LC_10_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4604\,
            lcout => \o_X_c_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_1__nesr_4C_net\,
            ce => \N__6575\,
            sr => \N__6511\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_0_0_c_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4865\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_17_0_\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_1_0_c_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4874\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_0\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_2_0_c_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4892\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_1\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_549\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_549_THRU_LUT4_0_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4883\,
            in3 => \N__4232\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_549_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_549\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_550\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_550_THRU_LUT4_0_LC_11_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4829\,
            in3 => \N__4391\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_550_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_550\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_4_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_4_0_c_RNIQ3MM_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5018\,
            in3 => \N__4379\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_551\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_4_6\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_5_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_5_0_c_RNIGV3E_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4835\,
            in2 => \N__4844\,
            in3 => \N__4364\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_552\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_5_6\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_553\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_553_THRU_LUT4_0_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5027\,
            in3 => \N__4352\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_553_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_553\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_554\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_554_THRU_LUT4_0_LC_11_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5036\,
            in3 => \N__4343\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_554_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_11_18_0_\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_555\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_555_THRU_LUT4_0_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5105\,
            in3 => \N__4331\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_555_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_555\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_556\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_556_THRU_LUT4_0_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5009\,
            in3 => \N__4316\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_556_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_556\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_557\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_557_THRU_LUT4_0_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5360\,
            in3 => \N__4301\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_557_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_557\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_558\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_558_THRU_LUT4_0_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5522\,
            in2 => \_gnd_net_\,
            in3 => \N__4505\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_558_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_558\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_559\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_559_THRU_LUT4_0_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4529\,
            in2 => \_gnd_net_\,
            in3 => \N__4493\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_559_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_559\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_560\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_11_0_c_RNIHNIP_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4490\,
            in2 => \_gnd_net_\,
            in3 => \N__4484\,
            lcout => \DFT.multiplier.regsA_un3_result_axb_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_0_0_c_RNO_LC_11_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5868\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5246\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_655\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_655_THRU_LUT4_0_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5291\,
            in3 => \N__4448\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_655_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_655\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_656\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_656_THRU_LUT4_0_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5282\,
            in3 => \N__4436\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_656_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_656\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_657\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_657_THRU_LUT4_0_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5264\,
            in3 => \N__4421\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_657_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_657\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_658\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_658_THRU_LUT4_0_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5255\,
            in3 => \N__4406\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_658_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_658\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_4_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_4_0_c_RNIICTH_LC_11_19_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4991\,
            in2 => \N__5273\,
            in3 => \N__4571\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_659\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_4_7\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_5_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_5_0_c_RNIUORI_LC_11_19_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5297\,
            in2 => \_gnd_net_\,
            in3 => \N__4556\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_660\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_5_7\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_661\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_661_THRU_LUT4_0_LC_11_19_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5498\,
            in2 => \_gnd_net_\,
            in3 => \N__4544\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_661_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_661\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_662\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_662_THRU_LUT4_0_LC_11_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4541\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_662_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_13_0_c_RNO_LC_11_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5944\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_13_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.state_RNIR1CE_0_LC_11_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5166\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5207\,
            lcout => \DFT.state_2_0\,
            ltout => \DFT.state_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.state_RNITIC91_1_LC_11_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__6530\,
            in1 => \N__5167\,
            in2 => \N__4520\,
            in3 => \N__5065\,
            lcout => \DFT.un1_state_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.state_0_LC_11_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5091\,
            lcout => \DFT.stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.state_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.state_1_LC_11_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__5092\,
            in1 => \N__5165\,
            in2 => \_gnd_net_\,
            in3 => \N__5066\,
            lcout => \DFT.stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.state_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_11_0_c_RNO_LC_11_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5943\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.o_X_0__nesr_7_LC_11_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4657\,
            lcout => \X_0__7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_0__nesr_7C_net\,
            ce => \N__5632\,
            sr => \N__6497\
        );

    \DFT.o_X_0__nesr_9_LC_11_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4645\,
            lcout => \X_0__9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_0__nesr_7C_net\,
            ce => \N__5632\,
            sr => \N__6497\
        );

    \DFT.o_X_0__nesr_8_LC_11_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4634\,
            lcout => \X_0__8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_0__nesr_7C_net\,
            ce => \N__5632\,
            sr => \N__6497\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_RNIRG904_LC_11_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5237\,
            in2 => \N__5456\,
            in3 => \N__4789\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNIRG904\,
            ltout => OPEN,
            carryin => \bfn_11_22_0_\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.regsA_un3_result_cry_2_THRU_LUT4_0_LC_11_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4622\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.o_X_1__nesr_10_LC_11_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6143\,
            in2 => \N__5341\,
            in3 => \_gnd_net_\,
            lcout => \X_1__10\,
            ltout => OPEN,
            carryin => \bfn_11_23_0_\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_2_0\,
            clk => \INVDFT.o_X_1__nesr_10C_net\,
            ce => \N__4762\,
            sr => \N__6504\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_2_c_RNI1KHL1_LC_11_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6104\,
            in2 => \N__4592\,
            in3 => \N__4583\,
            lcout => \DFT.x_11\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_2_0\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIGSDC2_LC_11_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5489\,
            in2 => \N__4820\,
            in3 => \N__4811\,
            lcout => \DFT.x_12\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_3\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_4_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNI7QS33_LC_11_23_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5474\,
            in2 => \N__4808\,
            in3 => \N__4799\,
            lcout => \DFT.x_13\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_4_0\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_5_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIEKOF6_LC_11_23_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4796\,
            in2 => \N__4790\,
            in3 => \N__4775\,
            lcout => \DFT.x_14\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_5_0\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_6_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNIS7913_LC_11_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4772\,
            in2 => \_gnd_net_\,
            in3 => \N__4766\,
            lcout => \DFT.x_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.o_X_1__nesr_15_LC_11_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4681\,
            lcout => \X_1__15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_1__nesr_10C_net\,
            ce => \N__4762\,
            sr => \N__6504\
        );

    \DFT.o_X_1__nesr_14_LC_11_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5323\,
            lcout => \X_1__14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_1__nesr_10C_net\,
            ce => \N__4762\,
            sr => \N__6504\
        );

    \DFT.o_X_0__nesr_13_LC_11_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4705\,
            lcout => \X_0__13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_0__nesr_13C_net\,
            ce => \N__5639\,
            sr => \N__6508\
        );

    \DFT.o_X_0__nesr_12_LC_11_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4693\,
            lcout => \X_0__12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_0__nesr_13C_net\,
            ce => \N__5639\,
            sr => \N__6508\
        );

    \DFT.o_X_0__nesr_15_LC_11_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4682\,
            lcout => \X_0__15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_0__nesr_13C_net\,
            ce => \N__5639\,
            sr => \N__6508\
        );

    \o_X_0__nesr_9_LC_11_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4985\,
            lcout => \o_X_c_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_0__nesr_9C_net\,
            ce => \N__6576\,
            sr => \N__6513\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_2_0_c_RNO_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5835\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_3_0_c_RNO_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5836\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_1_0_c_RNO_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5834\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_0_0_c_RNO_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5833\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_4_0_c_RNO_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_6_b_l_ofx_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6032\,
            in3 => \N__5839\,
            lcout => \DFT.multiplier.regsA_un3_result_6_b_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_6_ma_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5840\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_6_ma_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_4_0_c_RNO_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5838\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.b_6_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000101011101010"
        )
    port map (
            in0 => \N__6014\,
            in1 => \N__5221\,
            in2 => \N__5171\,
            in3 => \N__5077\,
            lcout => \DFT.bZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.b_6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_9_0_c_RNO_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5876\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.a_0_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__5879\,
            in1 => \N__5096\,
            in2 => \_gnd_net_\,
            in3 => \N__5076\,
            lcout => \DFT.aZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.b_6C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_8_0_c_RNO_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5875\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_7_0_c_RNO_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5874\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_5_ma_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5873\,
            in2 => \_gnd_net_\,
            in3 => \N__6013\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_5_ma_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_10_0_c_RNO_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5877\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_10_0_c_RNO_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5878\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_5_b_l_ofx_LC_12_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5885\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6026\,
            lcout => \DFT.multiplier.regsA_un3_result_5_b_l_ofx_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_6_ma_LC_12_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6027\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5887\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_6_ma_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_1_0_c_RNO_LC_12_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5881\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_2_0_c_RNO_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5882\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_5_ma_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5886\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_5_ma_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_3_0_c_RNO_LC_12_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5883\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_4_0_c_RNO_LC_12_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5884\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_RNO_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5880\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5366\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_763\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_763_THRU_LUT4_0_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5348\,
            in2 => \_gnd_net_\,
            in3 => \N__5225\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_763_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_763\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_764\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_1_0_c_RNIV67N_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__5423\,
            in1 => \N__5951\,
            in2 => \N__5954\,
            in3 => \N__5381\,
            lcout => \DFT.multiplier.regsA_un3_result_axb_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_RNO_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5946\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_11_0_c_RNO_LC_12_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5945\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_1_0_c_RNO_LC_12_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5947\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.o_X_0__nesr_10_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6142\,
            in2 => \_gnd_net_\,
            in3 => \N__5342\,
            lcout => \X_0__10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_0__nesr_10C_net\,
            ce => \N__5634\,
            sr => \N__6505\
        );

    \DFT.o_X_0__nesr_14_LC_12_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5324\,
            lcout => \X_0__14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_0__nesr_14C_net\,
            ce => \N__5633\,
            sr => \N__6509\
        );

    \DFT.o_X_0__nesr_11_LC_12_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5308\,
            lcout => \X_0__11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_0__nesr_11C_net\,
            ce => \N__5638\,
            sr => \N__6512\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_6_a_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5942\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6035\,
            lcout => \DFT.multiplier.regsA_un3_result_6_a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_3_0_c_RNO_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5941\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_RNILH0D_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5531\,
            in2 => \N__6077\,
            in3 => \N__6076\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_897\,
            ltout => OPEN,
            carryin => \bfn_13_17_0_\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_2_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_2_c_RNII9QL_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6053\,
            in2 => \N__6206\,
            in3 => \N__5459\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_898\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_2_2\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_3_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_3_c_RNIR3291_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6389\,
            in2 => \N__6188\,
            in3 => \N__5438\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_899\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_3_1\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_4_c_RNI9M7E_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110100110010110"
        )
    port map (
            in0 => \N__6170\,
            in1 => \N__6377\,
            in2 => \N__5435\,
            in3 => \N__5426\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_900\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_RNO_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5870\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_7_0_c_RNO_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5872\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_5_b_l_ofx_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5869\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6018\,
            lcout => \DFT.multiplier.regsA_un3_result_5_b_l_ofx_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_6_ma_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6033\,
            in3 => \N__5871\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_6_ma_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_1_0_c_RNO_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5889\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_3_0_c_RNO_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5893\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_5_b_l_ofx_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6028\,
            in2 => \_gnd_net_\,
            in3 => \N__5895\,
            lcout => \DFT.multiplier.regsA_un3_result_5_b_l_ofx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_1_0_c_RNO_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5890\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_0_0_c_RNO_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5888\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_2_0_c_RNO_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5892\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_4_0_c_RNO_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5894\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_2_0_c_RNO_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5891\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_12_0_c_RNO_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5902\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_12_0_c_RNO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_9_0_c_RNO_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5899\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_7_0_c_RNO_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5900\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_5_b_l_ofx_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5896\,
            in2 => \_gnd_net_\,
            in3 => \N__6022\,
            lcout => \DFT.multiplier.regsA_un3_result_5_b_l_ofx_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_6_ma_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__5897\,
            in1 => \_gnd_net_\,
            in2 => \N__6034\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_6_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_5_ma_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5901\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_5_ma\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_8_0_c_RNO_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__5898\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.o_X_0__nesr_6_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5687\,
            in2 => \_gnd_net_\,
            in3 => \N__5663\,
            lcout => \X_0__6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVDFT.o_X_0__nesr_6C_net\,
            ce => \N__5622\,
            sr => \N__6500\
        );

    \o_X_0__nesr_7_LC_13_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5582\,
            lcout => \o_X_c_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_0__nesr_7C_net\,
            ce => \N__6580\,
            sr => \N__6517\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5549\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_17_0_\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_727\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_727_THRU_LUT4_0_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5540\,
            in3 => \N__5525\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_727_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_727\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_728\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_728_THRU_LUT4_0_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6212\,
            in2 => \_gnd_net_\,
            in3 => \N__6197\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_728_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_728\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_729\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_729_THRU_LUT4_0_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6194\,
            in2 => \_gnd_net_\,
            in3 => \N__6176\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_729_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_729\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_730\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_730_THRU_LUT4_0_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6173\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_730_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_0_0_c_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6161\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_14_18_0_\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_691\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_LUT4_0_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6152\,
            in3 => \N__6116\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_691\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_692\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_692_THRU_LUT4_0_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6113\,
            in3 => \N__6089\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_692_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_692\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_693\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_LUT4_0_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6086\,
            in3 => \N__6062\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_693\,
            carryout => \DFT.multiplier.mult1_AdderTree2i_bigtree_694\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.mult1_AdderTree2i_bigtree_694_THRU_LUT4_0_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6059\,
            in2 => \_gnd_net_\,
            in3 => \N__6047\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_694_THRU_CO\,
            ltout => OPEN,
            carryin => \DFT.multiplier.mult1_AdderTree2i_bigtree_694\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_4_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_4_0_c_RNIJ7TP_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6404\,
            in2 => \N__6398\,
            in3 => \N__6383\,
            lcout => \DFT.multiplier.mult1_AdderTree2i_bigtree_695\,
            ltout => OPEN,
            carryin => \DFT.multiplier.regsA_un3_result_cry_4_3\,
            carryout => \DFT.multiplier.regsA_un3_result_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DFT.multiplier.regsA_un3_result_cry_5_THRU_LUT4_0_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6380\,
            lcout => \DFT.multiplier.regsA_un3_result_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \o_X_0__nesr_1_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6371\,
            lcout => \o_X_c_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_0__nesr_1C_net\,
            ce => \N__6570\,
            sr => \N__6501\
        );

    \o_X_0__nesr_0_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6338\,
            lcout => \o_X_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_0__nesr_1C_net\,
            ce => \N__6570\,
            sr => \N__6501\
        );

    \o_X_1__nesr_8_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6311\,
            lcout => \o_X_c_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_1__nesr_8C_net\,
            ce => \N__6572\,
            sr => \N__6506\
        );

    \o_X_0__nesr_3_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6278\,
            lcout => \o_X_c_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_0__nesr_3C_net\,
            ce => \N__6574\,
            sr => \N__6510\
        );

    \o_X_0__nesr_2_LC_14_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6257\,
            lcout => \o_X_c_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_0__nesr_3C_net\,
            ce => \N__6574\,
            sr => \N__6510\
        );

    \o_X_0__nesr_4_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6236\,
            lcout => \o_X_c_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_0__nesr_4C_net\,
            ce => \N__6577\,
            sr => \N__6514\
        );

    \o_X_0__nesr_8_LC_14_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6743\,
            lcout => \o_X_c_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_0__nesr_8C_net\,
            ce => \N__6579\,
            sr => \N__6516\
        );

    \o_X_1__nesr_9_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6710\,
            lcout => \o_X_c_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_1__nesr_9C_net\,
            ce => \N__6578\,
            sr => \N__6515\
        );

    \o_X_0__nesr_5_LC_15_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6629\,
            lcout => \o_X_c_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_0__nesr_5C_net\,
            ce => \N__6581\,
            sr => \N__6518\
        );

    \o_X_0__nesr_6_LC_15_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__6605\,
            lcout => \o_X_c_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVo_X_0__nesr_5C_net\,
            ce => \N__6581\,
            sr => \N__6518\
        );

    \CONSTANT_ONE_LUT4_LC_16_32_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
