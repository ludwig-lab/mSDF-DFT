// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 12 2024 10:20:51

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "top_test" view "INTERFACE"

module top_test (
    o_X,
    i_ref_clk,
    done,
    i_rst);

    output [31:0] o_X;
    input i_ref_clk;
    output done;
    input i_rst;

    wire N__7068;
    wire N__7067;
    wire N__7066;
    wire N__7059;
    wire N__7058;
    wire N__7057;
    wire N__7050;
    wire N__7049;
    wire N__7048;
    wire N__7041;
    wire N__7040;
    wire N__7039;
    wire N__7032;
    wire N__7031;
    wire N__7030;
    wire N__7023;
    wire N__7022;
    wire N__7021;
    wire N__7014;
    wire N__7013;
    wire N__7012;
    wire N__7005;
    wire N__7004;
    wire N__7003;
    wire N__6996;
    wire N__6995;
    wire N__6994;
    wire N__6987;
    wire N__6986;
    wire N__6985;
    wire N__6978;
    wire N__6977;
    wire N__6976;
    wire N__6969;
    wire N__6968;
    wire N__6967;
    wire N__6960;
    wire N__6959;
    wire N__6958;
    wire N__6951;
    wire N__6950;
    wire N__6949;
    wire N__6942;
    wire N__6941;
    wire N__6940;
    wire N__6933;
    wire N__6932;
    wire N__6931;
    wire N__6924;
    wire N__6923;
    wire N__6922;
    wire N__6915;
    wire N__6914;
    wire N__6913;
    wire N__6906;
    wire N__6905;
    wire N__6904;
    wire N__6897;
    wire N__6896;
    wire N__6895;
    wire N__6888;
    wire N__6887;
    wire N__6886;
    wire N__6879;
    wire N__6878;
    wire N__6877;
    wire N__6870;
    wire N__6869;
    wire N__6868;
    wire N__6861;
    wire N__6860;
    wire N__6859;
    wire N__6852;
    wire N__6851;
    wire N__6850;
    wire N__6843;
    wire N__6842;
    wire N__6841;
    wire N__6834;
    wire N__6833;
    wire N__6832;
    wire N__6825;
    wire N__6824;
    wire N__6823;
    wire N__6816;
    wire N__6815;
    wire N__6814;
    wire N__6807;
    wire N__6806;
    wire N__6805;
    wire N__6798;
    wire N__6797;
    wire N__6796;
    wire N__6789;
    wire N__6788;
    wire N__6787;
    wire N__6780;
    wire N__6779;
    wire N__6778;
    wire N__6771;
    wire N__6770;
    wire N__6769;
    wire N__6762;
    wire N__6761;
    wire N__6760;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6734;
    wire N__6731;
    wire N__6728;
    wire N__6725;
    wire N__6722;
    wire N__6719;
    wire N__6716;
    wire N__6713;
    wire N__6710;
    wire N__6707;
    wire N__6704;
    wire N__6701;
    wire N__6698;
    wire N__6697;
    wire N__6696;
    wire N__6695;
    wire N__6692;
    wire N__6689;
    wire N__6686;
    wire N__6685;
    wire N__6684;
    wire N__6683;
    wire N__6680;
    wire N__6673;
    wire N__6670;
    wire N__6667;
    wire N__6664;
    wire N__6661;
    wire N__6652;
    wire N__6649;
    wire N__6646;
    wire N__6641;
    wire N__6638;
    wire N__6635;
    wire N__6632;
    wire N__6629;
    wire N__6626;
    wire N__6623;
    wire N__6620;
    wire N__6617;
    wire N__6614;
    wire N__6611;
    wire N__6608;
    wire N__6605;
    wire N__6602;
    wire N__6599;
    wire N__6596;
    wire N__6593;
    wire N__6590;
    wire N__6587;
    wire N__6584;
    wire N__6581;
    wire N__6580;
    wire N__6579;
    wire N__6578;
    wire N__6577;
    wire N__6576;
    wire N__6575;
    wire N__6574;
    wire N__6573;
    wire N__6572;
    wire N__6571;
    wire N__6570;
    wire N__6569;
    wire N__6568;
    wire N__6567;
    wire N__6536;
    wire N__6533;
    wire N__6530;
    wire N__6529;
    wire N__6528;
    wire N__6525;
    wire N__6522;
    wire N__6519;
    wire N__6518;
    wire N__6517;
    wire N__6516;
    wire N__6515;
    wire N__6514;
    wire N__6513;
    wire N__6512;
    wire N__6511;
    wire N__6510;
    wire N__6509;
    wire N__6508;
    wire N__6507;
    wire N__6506;
    wire N__6505;
    wire N__6504;
    wire N__6503;
    wire N__6502;
    wire N__6501;
    wire N__6500;
    wire N__6499;
    wire N__6498;
    wire N__6497;
    wire N__6496;
    wire N__6495;
    wire N__6492;
    wire N__6491;
    wire N__6490;
    wire N__6487;
    wire N__6484;
    wire N__6425;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6371;
    wire N__6368;
    wire N__6365;
    wire N__6362;
    wire N__6359;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6344;
    wire N__6341;
    wire N__6338;
    wire N__6335;
    wire N__6332;
    wire N__6329;
    wire N__6326;
    wire N__6323;
    wire N__6320;
    wire N__6317;
    wire N__6314;
    wire N__6311;
    wire N__6308;
    wire N__6305;
    wire N__6302;
    wire N__6299;
    wire N__6296;
    wire N__6293;
    wire N__6290;
    wire N__6287;
    wire N__6284;
    wire N__6281;
    wire N__6278;
    wire N__6275;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6263;
    wire N__6260;
    wire N__6257;
    wire N__6254;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6242;
    wire N__6239;
    wire N__6236;
    wire N__6233;
    wire N__6230;
    wire N__6227;
    wire N__6224;
    wire N__6221;
    wire N__6218;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6203;
    wire N__6200;
    wire N__6197;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6182;
    wire N__6179;
    wire N__6176;
    wire N__6173;
    wire N__6170;
    wire N__6167;
    wire N__6164;
    wire N__6161;
    wire N__6158;
    wire N__6155;
    wire N__6152;
    wire N__6149;
    wire N__6146;
    wire N__6143;
    wire N__6142;
    wire N__6139;
    wire N__6136;
    wire N__6133;
    wire N__6130;
    wire N__6127;
    wire N__6124;
    wire N__6121;
    wire N__6116;
    wire N__6113;
    wire N__6110;
    wire N__6107;
    wire N__6104;
    wire N__6101;
    wire N__6098;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6077;
    wire N__6076;
    wire N__6073;
    wire N__6070;
    wire N__6067;
    wire N__6062;
    wire N__6059;
    wire N__6056;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6041;
    wire N__6038;
    wire N__6035;
    wire N__6034;
    wire N__6033;
    wire N__6032;
    wire N__6029;
    wire N__6028;
    wire N__6027;
    wire N__6026;
    wire N__6023;
    wire N__6022;
    wire N__6019;
    wire N__6018;
    wire N__6015;
    wire N__6014;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6002;
    wire N__5997;
    wire N__5992;
    wire N__5989;
    wire N__5984;
    wire N__5969;
    wire N__5966;
    wire N__5963;
    wire N__5960;
    wire N__5957;
    wire N__5954;
    wire N__5953;
    wire N__5952;
    wire N__5951;
    wire N__5948;
    wire N__5947;
    wire N__5946;
    wire N__5945;
    wire N__5944;
    wire N__5943;
    wire N__5942;
    wire N__5941;
    wire N__5936;
    wire N__5935;
    wire N__5934;
    wire N__5933;
    wire N__5932;
    wire N__5931;
    wire N__5930;
    wire N__5929;
    wire N__5928;
    wire N__5927;
    wire N__5926;
    wire N__5925;
    wire N__5922;
    wire N__5913;
    wire N__5908;
    wire N__5903;
    wire N__5902;
    wire N__5901;
    wire N__5900;
    wire N__5899;
    wire N__5898;
    wire N__5897;
    wire N__5896;
    wire N__5895;
    wire N__5894;
    wire N__5893;
    wire N__5892;
    wire N__5891;
    wire N__5890;
    wire N__5889;
    wire N__5888;
    wire N__5887;
    wire N__5886;
    wire N__5885;
    wire N__5884;
    wire N__5883;
    wire N__5882;
    wire N__5881;
    wire N__5880;
    wire N__5879;
    wire N__5878;
    wire N__5877;
    wire N__5876;
    wire N__5875;
    wire N__5874;
    wire N__5873;
    wire N__5872;
    wire N__5871;
    wire N__5870;
    wire N__5869;
    wire N__5868;
    wire N__5865;
    wire N__5848;
    wire N__5841;
    wire N__5840;
    wire N__5839;
    wire N__5838;
    wire N__5837;
    wire N__5836;
    wire N__5835;
    wire N__5834;
    wire N__5833;
    wire N__5826;
    wire N__5823;
    wire N__5808;
    wire N__5791;
    wire N__5774;
    wire N__5759;
    wire N__5750;
    wire N__5747;
    wire N__5740;
    wire N__5723;
    wire N__5702;
    wire N__5699;
    wire N__5696;
    wire N__5693;
    wire N__5690;
    wire N__5687;
    wire N__5686;
    wire N__5683;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5663;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5650;
    wire N__5647;
    wire N__5644;
    wire N__5639;
    wire N__5638;
    wire N__5635;
    wire N__5634;
    wire N__5633;
    wire N__5632;
    wire N__5629;
    wire N__5626;
    wire N__5623;
    wire N__5622;
    wire N__5619;
    wire N__5616;
    wire N__5609;
    wire N__5606;
    wire N__5601;
    wire N__5596;
    wire N__5593;
    wire N__5590;
    wire N__5587;
    wire N__5582;
    wire N__5579;
    wire N__5576;
    wire N__5573;
    wire N__5570;
    wire N__5567;
    wire N__5564;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5552;
    wire N__5549;
    wire N__5546;
    wire N__5543;
    wire N__5540;
    wire N__5537;
    wire N__5534;
    wire N__5531;
    wire N__5528;
    wire N__5525;
    wire N__5522;
    wire N__5519;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5498;
    wire N__5495;
    wire N__5492;
    wire N__5489;
    wire N__5486;
    wire N__5483;
    wire N__5480;
    wire N__5477;
    wire N__5474;
    wire N__5471;
    wire N__5468;
    wire N__5465;
    wire N__5462;
    wire N__5459;
    wire N__5456;
    wire N__5453;
    wire N__5450;
    wire N__5447;
    wire N__5444;
    wire N__5441;
    wire N__5438;
    wire N__5435;
    wire N__5432;
    wire N__5429;
    wire N__5426;
    wire N__5423;
    wire N__5420;
    wire N__5417;
    wire N__5414;
    wire N__5411;
    wire N__5408;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5396;
    wire N__5393;
    wire N__5390;
    wire N__5387;
    wire N__5384;
    wire N__5381;
    wire N__5378;
    wire N__5375;
    wire N__5372;
    wire N__5369;
    wire N__5366;
    wire N__5363;
    wire N__5360;
    wire N__5357;
    wire N__5354;
    wire N__5351;
    wire N__5348;
    wire N__5345;
    wire N__5342;
    wire N__5341;
    wire N__5338;
    wire N__5335;
    wire N__5332;
    wire N__5329;
    wire N__5324;
    wire N__5323;
    wire N__5320;
    wire N__5317;
    wire N__5312;
    wire N__5309;
    wire N__5308;
    wire N__5305;
    wire N__5302;
    wire N__5297;
    wire N__5294;
    wire N__5291;
    wire N__5288;
    wire N__5285;
    wire N__5282;
    wire N__5279;
    wire N__5276;
    wire N__5273;
    wire N__5270;
    wire N__5267;
    wire N__5264;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5252;
    wire N__5249;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5221;
    wire N__5218;
    wire N__5217;
    wire N__5214;
    wire N__5211;
    wire N__5208;
    wire N__5207;
    wire N__5204;
    wire N__5201;
    wire N__5198;
    wire N__5195;
    wire N__5186;
    wire N__5183;
    wire N__5180;
    wire N__5179;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5171;
    wire N__5168;
    wire N__5167;
    wire N__5166;
    wire N__5165;
    wire N__5160;
    wire N__5157;
    wire N__5154;
    wire N__5147;
    wire N__5144;
    wire N__5141;
    wire N__5138;
    wire N__5135;
    wire N__5130;
    wire N__5125;
    wire N__5122;
    wire N__5119;
    wire N__5116;
    wire N__5111;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5092;
    wire N__5091;
    wire N__5088;
    wire N__5083;
    wire N__5078;
    wire N__5077;
    wire N__5076;
    wire N__5073;
    wire N__5072;
    wire N__5067;
    wire N__5066;
    wire N__5065;
    wire N__5062;
    wire N__5059;
    wire N__5056;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5027;
    wire N__5024;
    wire N__5021;
    wire N__5018;
    wire N__5015;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__5000;
    wire N__4997;
    wire N__4994;
    wire N__4991;
    wire N__4988;
    wire N__4985;
    wire N__4982;
    wire N__4979;
    wire N__4976;
    wire N__4975;
    wire N__4972;
    wire N__4969;
    wire N__4968;
    wire N__4963;
    wire N__4960;
    wire N__4959;
    wire N__4958;
    wire N__4955;
    wire N__4952;
    wire N__4949;
    wire N__4946;
    wire N__4939;
    wire N__4938;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4905;
    wire N__4902;
    wire N__4897;
    wire N__4892;
    wire N__4889;
    wire N__4886;
    wire N__4883;
    wire N__4880;
    wire N__4877;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4835;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4814;
    wire N__4811;
    wire N__4808;
    wire N__4805;
    wire N__4802;
    wire N__4799;
    wire N__4796;
    wire N__4793;
    wire N__4790;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4780;
    wire N__4775;
    wire N__4772;
    wire N__4769;
    wire N__4766;
    wire N__4763;
    wire N__4762;
    wire N__4759;
    wire N__4758;
    wire N__4755;
    wire N__4752;
    wire N__4751;
    wire N__4750;
    wire N__4747;
    wire N__4744;
    wire N__4741;
    wire N__4738;
    wire N__4735;
    wire N__4732;
    wire N__4725;
    wire N__4722;
    wire N__4719;
    wire N__4716;
    wire N__4713;
    wire N__4706;
    wire N__4705;
    wire N__4702;
    wire N__4699;
    wire N__4694;
    wire N__4693;
    wire N__4690;
    wire N__4687;
    wire N__4682;
    wire N__4681;
    wire N__4678;
    wire N__4675;
    wire N__4670;
    wire N__4667;
    wire N__4664;
    wire N__4661;
    wire N__4658;
    wire N__4657;
    wire N__4654;
    wire N__4651;
    wire N__4646;
    wire N__4645;
    wire N__4642;
    wire N__4639;
    wire N__4634;
    wire N__4633;
    wire N__4630;
    wire N__4627;
    wire N__4622;
    wire N__4619;
    wire N__4616;
    wire N__4613;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4601;
    wire N__4598;
    wire N__4595;
    wire N__4592;
    wire N__4589;
    wire N__4586;
    wire N__4583;
    wire N__4580;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4565;
    wire N__4562;
    wire N__4559;
    wire N__4556;
    wire N__4553;
    wire N__4550;
    wire N__4547;
    wire N__4544;
    wire N__4541;
    wire N__4538;
    wire N__4535;
    wire N__4532;
    wire N__4529;
    wire N__4526;
    wire N__4523;
    wire N__4520;
    wire N__4517;
    wire N__4514;
    wire N__4511;
    wire N__4508;
    wire N__4505;
    wire N__4502;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4484;
    wire N__4481;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4466;
    wire N__4463;
    wire N__4462;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4445;
    wire N__4442;
    wire N__4439;
    wire N__4436;
    wire N__4433;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4403;
    wire N__4400;
    wire N__4397;
    wire N__4394;
    wire N__4391;
    wire N__4388;
    wire N__4385;
    wire N__4382;
    wire N__4379;
    wire N__4376;
    wire N__4373;
    wire N__4370;
    wire N__4367;
    wire N__4364;
    wire N__4361;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4349;
    wire N__4346;
    wire N__4343;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4307;
    wire N__4304;
    wire N__4301;
    wire N__4298;
    wire N__4295;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4271;
    wire N__4268;
    wire N__4265;
    wire N__4262;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4250;
    wire N__4247;
    wire N__4244;
    wire N__4241;
    wire N__4238;
    wire N__4235;
    wire N__4232;
    wire N__4229;
    wire N__4226;
    wire N__4223;
    wire N__4222;
    wire N__4219;
    wire N__4216;
    wire N__4213;
    wire N__4208;
    wire N__4205;
    wire N__4202;
    wire N__4199;
    wire N__4196;
    wire N__4193;
    wire N__4190;
    wire N__4187;
    wire N__4184;
    wire N__4181;
    wire N__4178;
    wire N__4175;
    wire N__4172;
    wire N__4169;
    wire N__4166;
    wire N__4163;
    wire N__4160;
    wire N__4157;
    wire N__4154;
    wire N__4151;
    wire N__4148;
    wire N__4145;
    wire N__4142;
    wire N__4139;
    wire N__4136;
    wire N__4133;
    wire N__4130;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4115;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4007;
    wire N__4004;
    wire N__4001;
    wire N__3998;
    wire N__3995;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3983;
    wire N__3980;
    wire N__3977;
    wire N__3974;
    wire N__3971;
    wire N__3968;
    wire N__3965;
    wire N__3962;
    wire N__3959;
    wire N__3956;
    wire N__3953;
    wire N__3950;
    wire N__3947;
    wire N__3944;
    wire N__3941;
    wire N__3938;
    wire N__3935;
    wire N__3932;
    wire N__3929;
    wire N__3926;
    wire N__3923;
    wire N__3920;
    wire N__3917;
    wire N__3914;
    wire N__3911;
    wire N__3908;
    wire N__3905;
    wire N__3902;
    wire N__3899;
    wire N__3896;
    wire N__3893;
    wire N__3890;
    wire N__3887;
    wire N__3884;
    wire N__3881;
    wire N__3878;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3854;
    wire N__3851;
    wire N__3848;
    wire N__3845;
    wire N__3842;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3824;
    wire N__3821;
    wire N__3818;
    wire N__3815;
    wire N__3812;
    wire N__3809;
    wire N__3806;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3788;
    wire N__3785;
    wire N__3782;
    wire N__3779;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3767;
    wire N__3764;
    wire N__3761;
    wire N__3758;
    wire N__3755;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3713;
    wire N__3710;
    wire N__3707;
    wire N__3704;
    wire N__3701;
    wire N__3698;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3683;
    wire N__3680;
    wire N__3677;
    wire N__3674;
    wire N__3671;
    wire N__3668;
    wire N__3665;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3647;
    wire N__3644;
    wire N__3641;
    wire N__3638;
    wire N__3635;
    wire N__3632;
    wire N__3629;
    wire N__3626;
    wire N__3623;
    wire N__3620;
    wire N__3617;
    wire N__3614;
    wire N__3611;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3596;
    wire N__3593;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3569;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3548;
    wire N__3545;
    wire N__3542;
    wire N__3539;
    wire N__3536;
    wire N__3533;
    wire N__3530;
    wire N__3527;
    wire N__3524;
    wire N__3521;
    wire N__3518;
    wire N__3515;
    wire N__3514;
    wire N__3511;
    wire N__3508;
    wire N__3505;
    wire N__3502;
    wire N__3501;
    wire N__3496;
    wire N__3493;
    wire N__3490;
    wire N__3485;
    wire N__3482;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3470;
    wire N__3467;
    wire N__3464;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3431;
    wire N__3428;
    wire N__3425;
    wire N__3422;
    wire N__3419;
    wire N__3416;
    wire N__3413;
    wire N__3410;
    wire N__3407;
    wire N__3404;
    wire N__3401;
    wire N__3398;
    wire N__3395;
    wire N__3392;
    wire N__3389;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3377;
    wire N__3374;
    wire N__3371;
    wire N__3368;
    wire N__3365;
    wire N__3364;
    wire N__3363;
    wire N__3362;
    wire N__3361;
    wire N__3360;
    wire N__3359;
    wire N__3358;
    wire N__3357;
    wire N__3356;
    wire N__3355;
    wire N__3354;
    wire N__3353;
    wire N__3352;
    wire N__3351;
    wire N__3350;
    wire N__3349;
    wire N__3348;
    wire N__3347;
    wire N__3346;
    wire N__3345;
    wire N__3344;
    wire N__3343;
    wire N__3342;
    wire N__3341;
    wire N__3340;
    wire N__3339;
    wire N__3338;
    wire N__3337;
    wire N__3278;
    wire N__3275;
    wire N__3272;
    wire N__3269;
    wire N__3266;
    wire sys_clk_g;
    wire sys_clk;
    wire GNDG0;
    wire i_ref_clk_c;
    wire VCCG0;
    wire i_rst_c_i;
    wire \DFT.done_c_0 ;
    wire \DFT.o_done_RNOZ0Z_0_cascade_ ;
    wire done_c;
    wire \INVDFT.o_doneC_net ;
    wire \DFT.state_RNIHM3GZ0Z_0 ;
    wire o_X_c_18;
    wire o_X_c_16;
    wire INVo_X_1__nesr_2C_net;
    wire o_X_c_19;
    wire INVo_X_1__nesr_3C_net;
    wire o_X_c_21;
    wire INVo_X_1__nesr_5C_net;
    wire \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_2 ;
    wire bfn_9_19_0_;
    wire \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_2 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_619 ;
    wire \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_1 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_620 ;
    wire \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_1 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_621 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_0 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_622 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_ma_0 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_4 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_4 ;
    wire \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_625 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_626 ;
    wire bfn_9_20_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_627 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_628 ;
    wire \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO ;
    wire \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO ;
    wire X_1__8;
    wire \INVDFT.o_X_1__nesr_8C_net ;
    wire X_1__9;
    wire \INVDFT.o_X_1__nesr_7C_net ;
    wire X_1__7;
    wire o_X_c_17;
    wire o_X_c_23;
    wire INVo_X_1__nesr_1C_net;
    wire bfn_10_17_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_583 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_584 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_585 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_586 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_ma_1 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_5 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_5 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_589 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_590 ;
    wire bfn_10_18_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_591 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_592 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_593 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_594 ;
    wire \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_2 ;
    wire \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_3 ;
    wire \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_2 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_583_THRU_CO ;
    wire bfn_10_19_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_584_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_2_4 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_585_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_3_3 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_586_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_2 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_587 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_3 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_588 ;
    wire \DFT.multiplier.regsA_un3_result_cry_6_1 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_589_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_7_1 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_590_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_8_1 ;
    wire \DFT.multiplier.regsA_un3_result_cry_9_0 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_591_THRU_CO ;
    wire bfn_10_20_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_592_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_10_0 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_593_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_11 ;
    wire \DFT.multiplier.regsA_un3_result_axb_9 ;
    wire \DFT.multiplier.regsA_un3_result_cry_12 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_621_THRU_CO ;
    wire bfn_10_21_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_622_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_2_3 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_623 ;
    wire \DFT.multiplier.regsA_un3_result_cry_3_2 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_624 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_1 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_625_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_2 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_626_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_6_0 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_627_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_7_0 ;
    wire \DFT.multiplier.regsA_un3_result_cry_8 ;
    wire \DFT.multiplier.regsA_un3_result_cry_8_THRU_CO ;
    wire X_1__6;
    wire bfn_10_22_0_;
    wire \INVDFT.o_X_1__nesr_6C_net ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_620_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_824 ;
    wire \DFT.multiplier.regsA_un3_result_cry_2_1 ;
    wire \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNI8J5C1 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_825 ;
    wire \DFT.multiplier.regsA_un3_result_cry_3_0 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_826 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_860 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_8 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_827 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_861 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_1 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_828 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_862 ;
    wire \DFT.multiplier.regsA_un3_result_cry_6 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_829 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_863 ;
    wire \DFT.multiplier.regsA_un3_result_cry_7 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_830 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_864 ;
    wire \DFT.multiplier.regsA_un3_result_cry_8_0 ;
    wire \DFT.multiplier.regsA_un3_result_cry_9 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_831 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_865 ;
    wire bfn_10_23_0_;
    wire \DFT.multiplier.regsA_un3_result_axb_11 ;
    wire \DFT.multiplier.regsA_un3_result_cry_10 ;
    wire X_1__11;
    wire X_1__13;
    wire \INVDFT.o_X_1__nesr_12C_net ;
    wire X_1__12;
    wire o_X_c_22;
    wire INVo_X_1__nesr_6C_net;
    wire o_X_c_20;
    wire INVo_X_1__nesr_4C_net;
    wire bfn_11_17_0_;
    wire \DFT.multiplier.regsA_un3_result_cry_0 ;
    wire \DFT.multiplier.regsA_un3_result_cry_1 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_549_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_549 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_550_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_550 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_551 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_6 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_552 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_6 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_553_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_553 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_554 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_554_THRU_CO ;
    wire bfn_11_18_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_555_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_555 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_556_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_556 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_557_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_557 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_558_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_558 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_559_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_559 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_594_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_560 ;
    wire \DFT.multiplier.regsA_un3_result_axb_13 ;
    wire \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_3 ;
    wire bfn_11_19_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_655_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_655 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_656_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_656 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_657_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_657 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_658_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_658 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_659 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_7 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_660 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_7 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_661_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_661 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_662 ;
    wire bfn_11_20_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_662_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_13_0_c_RNO ;
    wire \DFT.state_2_0_cascade_ ;
    wire \INVDFT.state_0C_net ;
    wire \DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO ;
    wire \DFT.x_7 ;
    wire \DFT.x_9 ;
    wire \DFT.x_8 ;
    wire \INVDFT.o_X_0__nesr_7C_net ;
    wire bfn_11_22_0_;
    wire \DFT.multiplier.regsA_un3_result_cry_2 ;
    wire \DFT.multiplier.regsA_un3_result_cry_2_THRU_CO ;
    wire X_1__10;
    wire bfn_11_23_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_964 ;
    wire \DFT.multiplier.regsA_un3_result_cry_2_0 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_965 ;
    wire \DFT.multiplier.regsA_un3_result_cry_3 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_966 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_0 ;
    wire \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNIRG904 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_967 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_0 ;
    wire \DFT.multiplier.regsA_un3_result_axb_7 ;
    wire \DFT.multiplier.regsA_un3_result_cry_6_2 ;
    wire \INVDFT.o_X_1__nesr_10C_net ;
    wire \DFT.un1_state_1_0 ;
    wire \DFT.x_13 ;
    wire \DFT.x_12 ;
    wire \DFT.x_15 ;
    wire \INVDFT.o_X_0__nesr_13C_net ;
    wire X_0__15;
    wire o_X_c_15;
    wire INVo_X_0__nesr_9C_net;
    wire \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_3 ;
    wire \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_3 ;
    wire \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_4 ;
    wire \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_4 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_1 ;
    wire \DFT.multiplier.regsA_un3_result_6_b_l_ofx ;
    wire \DFT.multiplier.regsA_un3_result_cry_6_ma_1 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_2 ;
    wire \DFT.stateZ0Z_0 ;
    wire i_rst_c;
    wire \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_1 ;
    wire \DFT.state_2_0 ;
    wire \DFT.stateZ0Z_1 ;
    wire \INVDFT.b_6C_net ;
    wire \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_1 ;
    wire \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_1 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_ma_2 ;
    wire \DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO_0 ;
    wire \DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO ;
    wire \DFT.multiplier.regsA_un3_result_5_b_l_ofx_2 ;
    wire \DFT.multiplier.regsA_un3_result_cry_6_ma_2 ;
    wire \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_5 ;
    wire \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_4 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_ma_3 ;
    wire \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_4 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_3 ;
    wire \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_5 ;
    wire bfn_12_20_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_763_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_763 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_764 ;
    wire \DFT.multiplier.regsA_un3_result_axb_3 ;
    wire \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO ;
    wire \DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO_0 ;
    wire \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_963 ;
    wire \INVDFT.o_X_0__nesr_10C_net ;
    wire \DFT.x_14 ;
    wire \INVDFT.o_X_0__nesr_14C_net ;
    wire \DFT.x_11 ;
    wire \INVDFT.o_X_0__nesr_11C_net ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_897 ;
    wire bfn_13_17_0_;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_898 ;
    wire \DFT.multiplier.regsA_un3_result_cry_2_2 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_899 ;
    wire \DFT.multiplier.regsA_un3_result_cry_3_1 ;
    wire \DFT.multiplier.regsA_un3_result_6_a ;
    wire \DFT.multiplier.regsA_un3_result_cry_4 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_900 ;
    wire \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_0 ;
    wire \DFT.multiplier.regsA_un3_result_5_b_l_ofx_1 ;
    wire \DFT.multiplier.regsA_un3_result_cry_6_ma_0 ;
    wire \DFT.multiplier.regsA_un3_result_cry_12_0_c_RNO ;
    wire \DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_0 ;
    wire \DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_2 ;
    wire \DFT.multiplier.regsA_un3_result_5_b_l_ofx_0 ;
    wire \DFT.bZ0Z_6 ;
    wire \DFT.multiplier.regsA_un3_result_cry_6_ma ;
    wire \DFT.aZ0Z_0 ;
    wire \DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_0 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_823 ;
    wire \INVDFT.o_X_0__nesr_6C_net ;
    wire \DFT.un1_state_4_0 ;
    wire X_0__13;
    wire o_X_c_7;
    wire INVo_X_0__nesr_7C_net;
    wire \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_0 ;
    wire bfn_14_17_0_;
    wire \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_0 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_727_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_727 ;
    wire \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_728_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_728 ;
    wire \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_729_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_729 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_730 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_730_THRU_CO ;
    wire \DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_1 ;
    wire bfn_14_18_0_;
    wire \DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_1 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_691 ;
    wire \DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_0 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_692_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_692 ;
    wire \DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_0 ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_693 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_694_THRU_CO ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_694 ;
    wire \DFT.multiplier.regsA_un3_result_5_b_l_ofx ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_ma ;
    wire \DFT.multiplier.mult1_AdderTree2i_bigtree_695 ;
    wire \DFT.multiplier.regsA_un3_result_cry_4_3 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5 ;
    wire \DFT.multiplier.regsA_un3_result_cry_5_THRU_CO ;
    wire X_0__7;
    wire o_X_c_1;
    wire X_0__6;
    wire o_X_c_0;
    wire INVo_X_0__nesr_1C_net;
    wire X_1__14;
    wire o_X_c_24;
    wire INVo_X_1__nesr_8C_net;
    wire X_0__9;
    wire o_X_c_3;
    wire X_0__8;
    wire o_X_c_2;
    wire INVo_X_0__nesr_3C_net;
    wire X_0__10;
    wire o_X_c_4;
    wire INVo_X_0__nesr_4C_net;
    wire X_0__14;
    wire o_X_c_8;
    wire INVo_X_0__nesr_8C_net;
    wire X_1__15;
    wire o_X_c_31;
    wire INVo_X_1__nesr_9C_net;
    wire X_0__11;
    wire o_X_c_5;
    wire X_0__12;
    wire o_X_c_6;
    wire INVo_X_0__nesr_5C_net;
    wire done_c_0_g;
    wire i_rst_c_i_g;
    wire CONSTANT_ONE_NET;
    wire _gnd_net_;

    defparam pll.DELAY_ADJUSTMENT_MODE_FEEDBACK="FIXED";
    defparam pll.TEST_MODE=1'b0;
    defparam pll.SHIFTREG_DIV_MODE=2'b00;
    defparam pll.PLLOUT_SELECT="GENCLK";
    defparam pll.FILTER_RANGE=3'b010;
    defparam pll.FEEDBACK_PATH="SIMPLE";
    defparam pll.FDA_RELATIVE=4'b0000;
    defparam pll.FDA_FEEDBACK=4'b0000;
    defparam pll.ENABLE_ICEGATE=1'b0;
    defparam pll.DIVR=4'b0100;
    defparam pll.DIVQ=3'b101;
    defparam pll.DIVF=7'b0101111;
    defparam pll.DELAY_ADJUSTMENT_MODE_RELATIVE="FIXED";
    SB_PLL40_CORE pll (
            .EXTFEEDBACK(),
            .LATCHINPUTVALUE(),
            .SCLK(),
            .SDO(),
            .LOCK(),
            .PLLOUTCORE(sys_clk),
            .REFERENCECLK(N__3401),
            .RESETB(N__6419),
            .BYPASS(GNDG0),
            .SDI(),
            .DYNAMICDELAY({GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0,GNDG0}),
            .PLLOUTGLOBAL());
    IO_PAD o_X_obuf_29_iopad (
            .OE(N__7068),
            .DIN(N__7067),
            .DOUT(N__7066),
            .PACKAGEPIN(o_X[29]));
    defparam o_X_obuf_29_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_29_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_29_preio (
            .PADOEN(N__7068),
            .PADOUT(N__7067),
            .PADIN(N__7066),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6695),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_9_iopad (
            .OE(N__7059),
            .DIN(N__7058),
            .DOUT(N__7057),
            .PACKAGEPIN(o_X[9]));
    defparam o_X_obuf_9_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_9_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_9_preio (
            .PADOEN(N__7059),
            .PADOUT(N__7058),
            .PADIN(N__7057),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4968),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_26_iopad (
            .OE(N__7050),
            .DIN(N__7049),
            .DOUT(N__7048),
            .PACKAGEPIN(o_X[26]));
    defparam o_X_obuf_26_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_26_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_26_preio (
            .PADOEN(N__7050),
            .PADOUT(N__7049),
            .PADIN(N__7048),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6684),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_ref_clk_ibuf_iopad (
            .OE(N__7041),
            .DIN(N__7040),
            .DOUT(N__7039),
            .PACKAGEPIN(i_ref_clk));
    defparam i_ref_clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_ref_clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_ref_clk_ibuf_preio (
            .PADOEN(N__7041),
            .PADOUT(N__7040),
            .PADIN(N__7039),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_ref_clk_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_31_iopad (
            .OE(N__7032),
            .DIN(N__7031),
            .DOUT(N__7030),
            .PACKAGEPIN(o_X[31]));
    defparam o_X_obuf_31_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_31_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_31_preio (
            .PADOEN(N__7032),
            .PADOUT(N__7031),
            .PADIN(N__7030),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6697),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_7_iopad (
            .OE(N__7023),
            .DIN(N__7022),
            .DOUT(N__7021),
            .PACKAGEPIN(o_X[7]));
    defparam o_X_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_7_preio (
            .PADOEN(N__7023),
            .PADOUT(N__7022),
            .PADIN(N__7021),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__5570),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_13_iopad (
            .OE(N__7014),
            .DIN(N__7013),
            .DOUT(N__7012),
            .PACKAGEPIN(o_X[13]));
    defparam o_X_obuf_13_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_13_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_13_preio (
            .PADOEN(N__7014),
            .PADOUT(N__7013),
            .PADIN(N__7012),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4938),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_2_iopad (
            .OE(N__7005),
            .DIN(N__7004),
            .DOUT(N__7003),
            .PACKAGEPIN(o_X[2]));
    defparam o_X_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_2_preio (
            .PADOEN(N__7005),
            .PADOUT(N__7004),
            .PADIN(N__7003),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6248),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_14_iopad (
            .OE(N__6996),
            .DIN(N__6995),
            .DOUT(N__6994),
            .PACKAGEPIN(o_X[14]));
    defparam o_X_obuf_14_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_14_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_14_preio (
            .PADOEN(N__6996),
            .PADOUT(N__6995),
            .PADIN(N__6994),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4958),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_24_iopad (
            .OE(N__6987),
            .DIN(N__6986),
            .DOUT(N__6985),
            .PACKAGEPIN(o_X[24]));
    defparam o_X_obuf_24_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_24_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_24_preio (
            .PADOEN(N__6987),
            .PADOUT(N__6986),
            .PADIN(N__6985),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6299),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD i_rst_ibuf_iopad (
            .OE(N__6978),
            .DIN(N__6977),
            .DOUT(N__6976),
            .PACKAGEPIN(i_rst));
    defparam i_rst_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam i_rst_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO i_rst_ibuf_preio (
            .PADOEN(N__6978),
            .PADOUT(N__6977),
            .PADIN(N__6976),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(i_rst_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_5_iopad (
            .OE(N__6969),
            .DIN(N__6968),
            .DOUT(N__6967),
            .PACKAGEPIN(o_X[5]));
    defparam o_X_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_5_preio (
            .PADOEN(N__6969),
            .PADOUT(N__6968),
            .PADIN(N__6967),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6620),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_11_iopad (
            .OE(N__6960),
            .DIN(N__6959),
            .DOUT(N__6958),
            .PACKAGEPIN(o_X[11]));
    defparam o_X_obuf_11_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_11_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_11_preio (
            .PADOEN(N__6960),
            .PADOUT(N__6959),
            .PADIN(N__6958),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4975),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_27_iopad (
            .OE(N__6951),
            .DIN(N__6950),
            .DOUT(N__6949),
            .PACKAGEPIN(o_X[27]));
    defparam o_X_obuf_27_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_27_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_27_preio (
            .PADOEN(N__6951),
            .PADOUT(N__6950),
            .PADIN(N__6949),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6683),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_0_iopad (
            .OE(N__6942),
            .DIN(N__6941),
            .DOUT(N__6940),
            .PACKAGEPIN(o_X[0]));
    defparam o_X_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_0_preio (
            .PADOEN(N__6942),
            .PADOUT(N__6941),
            .PADIN(N__6940),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6332),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_22_iopad (
            .OE(N__6933),
            .DIN(N__6932),
            .DOUT(N__6931),
            .PACKAGEPIN(o_X[22]));
    defparam o_X_obuf_22_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_22_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_22_preio (
            .PADOEN(N__6933),
            .PADOUT(N__6932),
            .PADIN(N__6931),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4274),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_19_iopad (
            .OE(N__6924),
            .DIN(N__6923),
            .DOUT(N__6922),
            .PACKAGEPIN(o_X[19]));
    defparam o_X_obuf_19_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_19_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_19_preio (
            .PADOEN(N__6924),
            .PADOUT(N__6923),
            .PADIN(N__6922),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3434),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_28_iopad (
            .OE(N__6915),
            .DIN(N__6914),
            .DOUT(N__6913),
            .PACKAGEPIN(o_X[28]));
    defparam o_X_obuf_28_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_28_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_28_preio (
            .PADOEN(N__6915),
            .PADOUT(N__6914),
            .PADIN(N__6913),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6696),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_30_iopad (
            .OE(N__6906),
            .DIN(N__6905),
            .DOUT(N__6904),
            .PACKAGEPIN(o_X[30]));
    defparam o_X_obuf_30_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_30_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_30_preio (
            .PADOEN(N__6906),
            .PADOUT(N__6905),
            .PADIN(N__6904),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6698),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_8_iopad (
            .OE(N__6897),
            .DIN(N__6896),
            .DOUT(N__6895),
            .PACKAGEPIN(o_X[8]));
    defparam o_X_obuf_8_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_8_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_8_preio (
            .PADOEN(N__6897),
            .PADOUT(N__6896),
            .PADIN(N__6895),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6731),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD done_obuf_iopad (
            .OE(N__6888),
            .DIN(N__6887),
            .DOUT(N__6886),
            .PACKAGEPIN(done));
    defparam done_obuf_preio.NEG_TRIGGER=1'b0;
    defparam done_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO done_obuf_preio (
            .PADOEN(N__6888),
            .PADOUT(N__6887),
            .PADIN(N__6886),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3527),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_12_iopad (
            .OE(N__6879),
            .DIN(N__6878),
            .DOUT(N__6877),
            .PACKAGEPIN(o_X[12]));
    defparam o_X_obuf_12_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_12_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_12_preio (
            .PADOEN(N__6879),
            .PADOUT(N__6878),
            .PADIN(N__6877),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4959),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_3_iopad (
            .OE(N__6870),
            .DIN(N__6869),
            .DOUT(N__6868),
            .PACKAGEPIN(o_X[3]));
    defparam o_X_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_3_preio (
            .PADOEN(N__6870),
            .PADOUT(N__6869),
            .PADIN(N__6868),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6269),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_17_iopad (
            .OE(N__6861),
            .DIN(N__6860),
            .DOUT(N__6859),
            .PACKAGEPIN(o_X[17]));
    defparam o_X_obuf_17_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_17_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_17_preio (
            .PADOEN(N__6861),
            .PADOUT(N__6860),
            .PADIN(N__6859),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3677),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_25_iopad (
            .OE(N__6852),
            .DIN(N__6851),
            .DOUT(N__6850),
            .PACKAGEPIN(o_X[25]));
    defparam o_X_obuf_25_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_25_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_25_preio (
            .PADOEN(N__6852),
            .PADOUT(N__6851),
            .PADIN(N__6850),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6685),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_20_iopad (
            .OE(N__6843),
            .DIN(N__6842),
            .DOUT(N__6841),
            .PACKAGEPIN(o_X[20]));
    defparam o_X_obuf_20_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_20_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_20_preio (
            .PADOEN(N__6843),
            .PADOUT(N__6842),
            .PADIN(N__6841),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4262),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_6_iopad (
            .OE(N__6834),
            .DIN(N__6833),
            .DOUT(N__6832),
            .PACKAGEPIN(o_X[6]));
    defparam o_X_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_6_preio (
            .PADOEN(N__6834),
            .PADOUT(N__6833),
            .PADIN(N__6832),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6596),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_10_iopad (
            .OE(N__6825),
            .DIN(N__6824),
            .DOUT(N__6823),
            .PACKAGEPIN(o_X[10]));
    defparam o_X_obuf_10_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_10_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_10_preio (
            .PADOEN(N__6825),
            .PADOUT(N__6824),
            .PADIN(N__6823),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4976),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_1_iopad (
            .OE(N__6816),
            .DIN(N__6815),
            .DOUT(N__6814),
            .PACKAGEPIN(o_X[1]));
    defparam o_X_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_1_preio (
            .PADOEN(N__6816),
            .PADOUT(N__6815),
            .PADIN(N__6814),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6359),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_15_iopad (
            .OE(N__6807),
            .DIN(N__6806),
            .DOUT(N__6805),
            .PACKAGEPIN(o_X[15]));
    defparam o_X_obuf_15_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_15_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_15_preio (
            .PADOEN(N__6807),
            .PADOUT(N__6806),
            .PADIN(N__6805),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__4937),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_23_iopad (
            .OE(N__6798),
            .DIN(N__6797),
            .DOUT(N__6796),
            .PACKAGEPIN(o_X[23]));
    defparam o_X_obuf_23_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_23_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_23_preio (
            .PADOEN(N__6798),
            .PADOUT(N__6797),
            .PADIN(N__6796),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3659),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_18_iopad (
            .OE(N__6789),
            .DIN(N__6788),
            .DOUT(N__6787),
            .PACKAGEPIN(o_X[18]));
    defparam o_X_obuf_18_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_18_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_18_preio (
            .PADOEN(N__6789),
            .PADOUT(N__6788),
            .PADIN(N__6787),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3470),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_4_iopad (
            .OE(N__6780),
            .DIN(N__6779),
            .DOUT(N__6778),
            .PACKAGEPIN(o_X[4]));
    defparam o_X_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_4_preio (
            .PADOEN(N__6780),
            .PADOUT(N__6779),
            .PADIN(N__6778),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6224),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_16_iopad (
            .OE(N__6771),
            .DIN(N__6770),
            .DOUT(N__6769),
            .PACKAGEPIN(o_X[16]));
    defparam o_X_obuf_16_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_16_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_16_preio (
            .PADOEN(N__6771),
            .PADOUT(N__6770),
            .PADIN(N__6769),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3452),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD o_X_obuf_21_iopad (
            .OE(N__6762),
            .DIN(N__6761),
            .DOUT(N__6760),
            .PACKAGEPIN(o_X[21]));
    defparam o_X_obuf_21_preio.NEG_TRIGGER=1'b0;
    defparam o_X_obuf_21_preio.PIN_TYPE=6'b011001;
    PRE_IO o_X_obuf_21_preio (
            .PADOEN(N__6762),
            .PADOUT(N__6761),
            .PADIN(N__6760),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3419),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__1467 (
            .O(N__6743),
            .I(N__6740));
    LocalMux I__1466 (
            .O(N__6740),
            .I(N__6737));
    Span4Mux_h I__1465 (
            .O(N__6737),
            .I(N__6734));
    Odrv4 I__1464 (
            .O(N__6734),
            .I(X_0__14));
    IoInMux I__1463 (
            .O(N__6731),
            .I(N__6728));
    LocalMux I__1462 (
            .O(N__6728),
            .I(N__6725));
    Span4Mux_s0_v I__1461 (
            .O(N__6725),
            .I(N__6722));
    Span4Mux_h I__1460 (
            .O(N__6722),
            .I(N__6719));
    Span4Mux_v I__1459 (
            .O(N__6719),
            .I(N__6716));
    Span4Mux_v I__1458 (
            .O(N__6716),
            .I(N__6713));
    Odrv4 I__1457 (
            .O(N__6713),
            .I(o_X_c_8));
    InMux I__1456 (
            .O(N__6710),
            .I(N__6707));
    LocalMux I__1455 (
            .O(N__6707),
            .I(N__6704));
    Span4Mux_h I__1454 (
            .O(N__6704),
            .I(N__6701));
    Odrv4 I__1453 (
            .O(N__6701),
            .I(X_1__15));
    IoInMux I__1452 (
            .O(N__6698),
            .I(N__6692));
    IoInMux I__1451 (
            .O(N__6697),
            .I(N__6689));
    IoInMux I__1450 (
            .O(N__6696),
            .I(N__6686));
    IoInMux I__1449 (
            .O(N__6695),
            .I(N__6680));
    LocalMux I__1448 (
            .O(N__6692),
            .I(N__6673));
    LocalMux I__1447 (
            .O(N__6689),
            .I(N__6673));
    LocalMux I__1446 (
            .O(N__6686),
            .I(N__6673));
    IoInMux I__1445 (
            .O(N__6685),
            .I(N__6670));
    IoInMux I__1444 (
            .O(N__6684),
            .I(N__6667));
    IoInMux I__1443 (
            .O(N__6683),
            .I(N__6664));
    LocalMux I__1442 (
            .O(N__6680),
            .I(N__6661));
    IoSpan4Mux I__1441 (
            .O(N__6673),
            .I(N__6652));
    LocalMux I__1440 (
            .O(N__6670),
            .I(N__6652));
    LocalMux I__1439 (
            .O(N__6667),
            .I(N__6652));
    LocalMux I__1438 (
            .O(N__6664),
            .I(N__6652));
    Span4Mux_s3_h I__1437 (
            .O(N__6661),
            .I(N__6649));
    IoSpan4Mux I__1436 (
            .O(N__6652),
            .I(N__6646));
    Span4Mux_v I__1435 (
            .O(N__6649),
            .I(N__6641));
    Span4Mux_s3_h I__1434 (
            .O(N__6646),
            .I(N__6641));
    Sp12to4 I__1433 (
            .O(N__6641),
            .I(N__6638));
    Span12Mux_h I__1432 (
            .O(N__6638),
            .I(N__6635));
    Span12Mux_v I__1431 (
            .O(N__6635),
            .I(N__6632));
    Odrv12 I__1430 (
            .O(N__6632),
            .I(o_X_c_31));
    InMux I__1429 (
            .O(N__6629),
            .I(N__6626));
    LocalMux I__1428 (
            .O(N__6626),
            .I(N__6623));
    Odrv12 I__1427 (
            .O(N__6623),
            .I(X_0__11));
    IoInMux I__1426 (
            .O(N__6620),
            .I(N__6617));
    LocalMux I__1425 (
            .O(N__6617),
            .I(N__6614));
    Sp12to4 I__1424 (
            .O(N__6614),
            .I(N__6611));
    Span12Mux_h I__1423 (
            .O(N__6611),
            .I(N__6608));
    Odrv12 I__1422 (
            .O(N__6608),
            .I(o_X_c_5));
    InMux I__1421 (
            .O(N__6605),
            .I(N__6602));
    LocalMux I__1420 (
            .O(N__6602),
            .I(N__6599));
    Odrv12 I__1419 (
            .O(N__6599),
            .I(X_0__12));
    IoInMux I__1418 (
            .O(N__6596),
            .I(N__6593));
    LocalMux I__1417 (
            .O(N__6593),
            .I(N__6590));
    Span12Mux_s5_h I__1416 (
            .O(N__6590),
            .I(N__6587));
    Span12Mux_h I__1415 (
            .O(N__6587),
            .I(N__6584));
    Odrv12 I__1414 (
            .O(N__6584),
            .I(o_X_c_6));
    CEMux I__1413 (
            .O(N__6581),
            .I(N__6536));
    CEMux I__1412 (
            .O(N__6580),
            .I(N__6536));
    CEMux I__1411 (
            .O(N__6579),
            .I(N__6536));
    CEMux I__1410 (
            .O(N__6578),
            .I(N__6536));
    CEMux I__1409 (
            .O(N__6577),
            .I(N__6536));
    CEMux I__1408 (
            .O(N__6576),
            .I(N__6536));
    CEMux I__1407 (
            .O(N__6575),
            .I(N__6536));
    CEMux I__1406 (
            .O(N__6574),
            .I(N__6536));
    CEMux I__1405 (
            .O(N__6573),
            .I(N__6536));
    CEMux I__1404 (
            .O(N__6572),
            .I(N__6536));
    CEMux I__1403 (
            .O(N__6571),
            .I(N__6536));
    CEMux I__1402 (
            .O(N__6570),
            .I(N__6536));
    CEMux I__1401 (
            .O(N__6569),
            .I(N__6536));
    CEMux I__1400 (
            .O(N__6568),
            .I(N__6536));
    CEMux I__1399 (
            .O(N__6567),
            .I(N__6536));
    GlobalMux I__1398 (
            .O(N__6536),
            .I(N__6533));
    gio2CtrlBuf I__1397 (
            .O(N__6533),
            .I(done_c_0_g));
    InMux I__1396 (
            .O(N__6530),
            .I(N__6525));
    InMux I__1395 (
            .O(N__6529),
            .I(N__6522));
    InMux I__1394 (
            .O(N__6528),
            .I(N__6519));
    LocalMux I__1393 (
            .O(N__6525),
            .I(N__6492));
    LocalMux I__1392 (
            .O(N__6522),
            .I(N__6487));
    LocalMux I__1391 (
            .O(N__6519),
            .I(N__6484));
    SRMux I__1390 (
            .O(N__6518),
            .I(N__6425));
    SRMux I__1389 (
            .O(N__6517),
            .I(N__6425));
    SRMux I__1388 (
            .O(N__6516),
            .I(N__6425));
    SRMux I__1387 (
            .O(N__6515),
            .I(N__6425));
    SRMux I__1386 (
            .O(N__6514),
            .I(N__6425));
    SRMux I__1385 (
            .O(N__6513),
            .I(N__6425));
    SRMux I__1384 (
            .O(N__6512),
            .I(N__6425));
    SRMux I__1383 (
            .O(N__6511),
            .I(N__6425));
    SRMux I__1382 (
            .O(N__6510),
            .I(N__6425));
    SRMux I__1381 (
            .O(N__6509),
            .I(N__6425));
    SRMux I__1380 (
            .O(N__6508),
            .I(N__6425));
    SRMux I__1379 (
            .O(N__6507),
            .I(N__6425));
    SRMux I__1378 (
            .O(N__6506),
            .I(N__6425));
    SRMux I__1377 (
            .O(N__6505),
            .I(N__6425));
    SRMux I__1376 (
            .O(N__6504),
            .I(N__6425));
    SRMux I__1375 (
            .O(N__6503),
            .I(N__6425));
    SRMux I__1374 (
            .O(N__6502),
            .I(N__6425));
    SRMux I__1373 (
            .O(N__6501),
            .I(N__6425));
    SRMux I__1372 (
            .O(N__6500),
            .I(N__6425));
    SRMux I__1371 (
            .O(N__6499),
            .I(N__6425));
    SRMux I__1370 (
            .O(N__6498),
            .I(N__6425));
    SRMux I__1369 (
            .O(N__6497),
            .I(N__6425));
    SRMux I__1368 (
            .O(N__6496),
            .I(N__6425));
    SRMux I__1367 (
            .O(N__6495),
            .I(N__6425));
    Glb2LocalMux I__1366 (
            .O(N__6492),
            .I(N__6425));
    SRMux I__1365 (
            .O(N__6491),
            .I(N__6425));
    SRMux I__1364 (
            .O(N__6490),
            .I(N__6425));
    Glb2LocalMux I__1363 (
            .O(N__6487),
            .I(N__6425));
    Glb2LocalMux I__1362 (
            .O(N__6484),
            .I(N__6425));
    GlobalMux I__1361 (
            .O(N__6425),
            .I(N__6422));
    gio2CtrlBuf I__1360 (
            .O(N__6422),
            .I(i_rst_c_i_g));
    IoInMux I__1359 (
            .O(N__6419),
            .I(N__6416));
    LocalMux I__1358 (
            .O(N__6416),
            .I(N__6413));
    IoSpan4Mux I__1357 (
            .O(N__6413),
            .I(N__6410));
    Span4Mux_s0_v I__1356 (
            .O(N__6410),
            .I(N__6407));
    Odrv4 I__1355 (
            .O(N__6407),
            .I(CONSTANT_ONE_NET));
    InMux I__1354 (
            .O(N__6404),
            .I(N__6401));
    LocalMux I__1353 (
            .O(N__6401),
            .I(\DFT.multiplier.regsA_un3_result_5_b_l_ofx ));
    CascadeMux I__1352 (
            .O(N__6398),
            .I(N__6395));
    InMux I__1351 (
            .O(N__6395),
            .I(N__6392));
    LocalMux I__1350 (
            .O(N__6392),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_ma ));
    InMux I__1349 (
            .O(N__6389),
            .I(N__6386));
    LocalMux I__1348 (
            .O(N__6386),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_695 ));
    InMux I__1347 (
            .O(N__6383),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_3 ));
    InMux I__1346 (
            .O(N__6380),
            .I(\DFT.multiplier.regsA_un3_result_cry_5 ));
    InMux I__1345 (
            .O(N__6377),
            .I(N__6374));
    LocalMux I__1344 (
            .O(N__6374),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_THRU_CO ));
    InMux I__1343 (
            .O(N__6371),
            .I(N__6368));
    LocalMux I__1342 (
            .O(N__6368),
            .I(N__6365));
    Span4Mux_h I__1341 (
            .O(N__6365),
            .I(N__6362));
    Odrv4 I__1340 (
            .O(N__6362),
            .I(X_0__7));
    IoInMux I__1339 (
            .O(N__6359),
            .I(N__6356));
    LocalMux I__1338 (
            .O(N__6356),
            .I(N__6353));
    IoSpan4Mux I__1337 (
            .O(N__6353),
            .I(N__6350));
    Span4Mux_s1_h I__1336 (
            .O(N__6350),
            .I(N__6347));
    Sp12to4 I__1335 (
            .O(N__6347),
            .I(N__6344));
    Span12Mux_h I__1334 (
            .O(N__6344),
            .I(N__6341));
    Odrv12 I__1333 (
            .O(N__6341),
            .I(o_X_c_1));
    InMux I__1332 (
            .O(N__6338),
            .I(N__6335));
    LocalMux I__1331 (
            .O(N__6335),
            .I(X_0__6));
    IoInMux I__1330 (
            .O(N__6332),
            .I(N__6329));
    LocalMux I__1329 (
            .O(N__6329),
            .I(N__6326));
    Span4Mux_s2_h I__1328 (
            .O(N__6326),
            .I(N__6323));
    Span4Mux_h I__1327 (
            .O(N__6323),
            .I(N__6320));
    Sp12to4 I__1326 (
            .O(N__6320),
            .I(N__6317));
    Span12Mux_v I__1325 (
            .O(N__6317),
            .I(N__6314));
    Odrv12 I__1324 (
            .O(N__6314),
            .I(o_X_c_0));
    InMux I__1323 (
            .O(N__6311),
            .I(N__6308));
    LocalMux I__1322 (
            .O(N__6308),
            .I(N__6305));
    Span4Mux_h I__1321 (
            .O(N__6305),
            .I(N__6302));
    Odrv4 I__1320 (
            .O(N__6302),
            .I(X_1__14));
    IoInMux I__1319 (
            .O(N__6299),
            .I(N__6296));
    LocalMux I__1318 (
            .O(N__6296),
            .I(N__6293));
    Span4Mux_s2_h I__1317 (
            .O(N__6293),
            .I(N__6290));
    Sp12to4 I__1316 (
            .O(N__6290),
            .I(N__6287));
    Span12Mux_v I__1315 (
            .O(N__6287),
            .I(N__6284));
    Span12Mux_h I__1314 (
            .O(N__6284),
            .I(N__6281));
    Odrv12 I__1313 (
            .O(N__6281),
            .I(o_X_c_24));
    InMux I__1312 (
            .O(N__6278),
            .I(N__6275));
    LocalMux I__1311 (
            .O(N__6275),
            .I(N__6272));
    Odrv4 I__1310 (
            .O(N__6272),
            .I(X_0__9));
    IoInMux I__1309 (
            .O(N__6269),
            .I(N__6266));
    LocalMux I__1308 (
            .O(N__6266),
            .I(N__6263));
    Span12Mux_s10_h I__1307 (
            .O(N__6263),
            .I(N__6260));
    Odrv12 I__1306 (
            .O(N__6260),
            .I(o_X_c_3));
    InMux I__1305 (
            .O(N__6257),
            .I(N__6254));
    LocalMux I__1304 (
            .O(N__6254),
            .I(N__6251));
    Odrv4 I__1303 (
            .O(N__6251),
            .I(X_0__8));
    IoInMux I__1302 (
            .O(N__6248),
            .I(N__6245));
    LocalMux I__1301 (
            .O(N__6245),
            .I(N__6242));
    Span12Mux_s9_h I__1300 (
            .O(N__6242),
            .I(N__6239));
    Odrv12 I__1299 (
            .O(N__6239),
            .I(o_X_c_2));
    InMux I__1298 (
            .O(N__6236),
            .I(N__6233));
    LocalMux I__1297 (
            .O(N__6233),
            .I(N__6230));
    Span4Mux_h I__1296 (
            .O(N__6230),
            .I(N__6227));
    Odrv4 I__1295 (
            .O(N__6227),
            .I(X_0__10));
    IoInMux I__1294 (
            .O(N__6224),
            .I(N__6221));
    LocalMux I__1293 (
            .O(N__6221),
            .I(N__6218));
    Span12Mux_s10_h I__1292 (
            .O(N__6218),
            .I(N__6215));
    Odrv12 I__1291 (
            .O(N__6215),
            .I(o_X_c_4));
    InMux I__1290 (
            .O(N__6212),
            .I(N__6209));
    LocalMux I__1289 (
            .O(N__6209),
            .I(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO ));
    CascadeMux I__1288 (
            .O(N__6206),
            .I(N__6203));
    InMux I__1287 (
            .O(N__6203),
            .I(N__6200));
    LocalMux I__1286 (
            .O(N__6200),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_728_THRU_CO ));
    InMux I__1285 (
            .O(N__6197),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_728 ));
    InMux I__1284 (
            .O(N__6194),
            .I(N__6191));
    LocalMux I__1283 (
            .O(N__6191),
            .I(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO ));
    CascadeMux I__1282 (
            .O(N__6188),
            .I(N__6185));
    InMux I__1281 (
            .O(N__6185),
            .I(N__6182));
    LocalMux I__1280 (
            .O(N__6182),
            .I(N__6179));
    Odrv4 I__1279 (
            .O(N__6179),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_729_THRU_CO ));
    InMux I__1278 (
            .O(N__6176),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_729 ));
    InMux I__1277 (
            .O(N__6173),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_730 ));
    InMux I__1276 (
            .O(N__6170),
            .I(N__6167));
    LocalMux I__1275 (
            .O(N__6167),
            .I(N__6164));
    Odrv4 I__1274 (
            .O(N__6164),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_730_THRU_CO ));
    CascadeMux I__1273 (
            .O(N__6161),
            .I(N__6158));
    InMux I__1272 (
            .O(N__6158),
            .I(N__6155));
    LocalMux I__1271 (
            .O(N__6155),
            .I(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_1 ));
    CascadeMux I__1270 (
            .O(N__6152),
            .I(N__6149));
    InMux I__1269 (
            .O(N__6149),
            .I(N__6146));
    LocalMux I__1268 (
            .O(N__6146),
            .I(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_1 ));
    InMux I__1267 (
            .O(N__6143),
            .I(N__6139));
    InMux I__1266 (
            .O(N__6142),
            .I(N__6136));
    LocalMux I__1265 (
            .O(N__6139),
            .I(N__6133));
    LocalMux I__1264 (
            .O(N__6136),
            .I(N__6130));
    Span4Mux_h I__1263 (
            .O(N__6133),
            .I(N__6127));
    Span4Mux_v I__1262 (
            .O(N__6130),
            .I(N__6124));
    Span4Mux_v I__1261 (
            .O(N__6127),
            .I(N__6121));
    Odrv4 I__1260 (
            .O(N__6124),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_CO ));
    Odrv4 I__1259 (
            .O(N__6121),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_CO ));
    InMux I__1258 (
            .O(N__6116),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_691 ));
    CascadeMux I__1257 (
            .O(N__6113),
            .I(N__6110));
    InMux I__1256 (
            .O(N__6110),
            .I(N__6107));
    LocalMux I__1255 (
            .O(N__6107),
            .I(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_0 ));
    InMux I__1254 (
            .O(N__6104),
            .I(N__6101));
    LocalMux I__1253 (
            .O(N__6101),
            .I(N__6098));
    Span4Mux_v I__1252 (
            .O(N__6098),
            .I(N__6095));
    Span4Mux_h I__1251 (
            .O(N__6095),
            .I(N__6092));
    Odrv4 I__1250 (
            .O(N__6092),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_692_THRU_CO ));
    InMux I__1249 (
            .O(N__6089),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_692 ));
    CascadeMux I__1248 (
            .O(N__6086),
            .I(N__6083));
    InMux I__1247 (
            .O(N__6083),
            .I(N__6080));
    LocalMux I__1246 (
            .O(N__6080),
            .I(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_0 ));
    CascadeMux I__1245 (
            .O(N__6077),
            .I(N__6073));
    InMux I__1244 (
            .O(N__6076),
            .I(N__6070));
    InMux I__1243 (
            .O(N__6073),
            .I(N__6067));
    LocalMux I__1242 (
            .O(N__6070),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_CO ));
    LocalMux I__1241 (
            .O(N__6067),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_CO ));
    InMux I__1240 (
            .O(N__6062),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_693 ));
    InMux I__1239 (
            .O(N__6059),
            .I(N__6056));
    LocalMux I__1238 (
            .O(N__6056),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO ));
    InMux I__1237 (
            .O(N__6053),
            .I(N__6050));
    LocalMux I__1236 (
            .O(N__6050),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_694_THRU_CO ));
    InMux I__1235 (
            .O(N__6047),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_694 ));
    InMux I__1234 (
            .O(N__6044),
            .I(N__6041));
    LocalMux I__1233 (
            .O(N__6041),
            .I(N__6038));
    Odrv12 I__1232 (
            .O(N__6038),
            .I(\DFT.multiplier.regsA_un3_result_5_b_l_ofx_0 ));
    InMux I__1231 (
            .O(N__6035),
            .I(N__6029));
    CascadeMux I__1230 (
            .O(N__6034),
            .I(N__6023));
    CascadeMux I__1229 (
            .O(N__6033),
            .I(N__6019));
    CascadeMux I__1228 (
            .O(N__6032),
            .I(N__6015));
    LocalMux I__1227 (
            .O(N__6029),
            .I(N__6010));
    InMux I__1226 (
            .O(N__6028),
            .I(N__6007));
    InMux I__1225 (
            .O(N__6027),
            .I(N__6002));
    InMux I__1224 (
            .O(N__6026),
            .I(N__6002));
    InMux I__1223 (
            .O(N__6023),
            .I(N__5997));
    InMux I__1222 (
            .O(N__6022),
            .I(N__5997));
    InMux I__1221 (
            .O(N__6019),
            .I(N__5992));
    InMux I__1220 (
            .O(N__6018),
            .I(N__5992));
    InMux I__1219 (
            .O(N__6015),
            .I(N__5989));
    InMux I__1218 (
            .O(N__6014),
            .I(N__5984));
    InMux I__1217 (
            .O(N__6013),
            .I(N__5984));
    Odrv4 I__1216 (
            .O(N__6010),
            .I(\DFT.bZ0Z_6 ));
    LocalMux I__1215 (
            .O(N__6007),
            .I(\DFT.bZ0Z_6 ));
    LocalMux I__1214 (
            .O(N__6002),
            .I(\DFT.bZ0Z_6 ));
    LocalMux I__1213 (
            .O(N__5997),
            .I(\DFT.bZ0Z_6 ));
    LocalMux I__1212 (
            .O(N__5992),
            .I(\DFT.bZ0Z_6 ));
    LocalMux I__1211 (
            .O(N__5989),
            .I(\DFT.bZ0Z_6 ));
    LocalMux I__1210 (
            .O(N__5984),
            .I(\DFT.bZ0Z_6 ));
    CascadeMux I__1209 (
            .O(N__5969),
            .I(N__5966));
    InMux I__1208 (
            .O(N__5966),
            .I(N__5963));
    LocalMux I__1207 (
            .O(N__5963),
            .I(N__5960));
    Span4Mux_h I__1206 (
            .O(N__5960),
            .I(N__5957));
    Odrv4 I__1205 (
            .O(N__5957),
            .I(\DFT.multiplier.regsA_un3_result_cry_6_ma ));
    CascadeMux I__1204 (
            .O(N__5954),
            .I(N__5948));
    InMux I__1203 (
            .O(N__5953),
            .I(N__5936));
    InMux I__1202 (
            .O(N__5952),
            .I(N__5936));
    InMux I__1201 (
            .O(N__5951),
            .I(N__5922));
    InMux I__1200 (
            .O(N__5948),
            .I(N__5913));
    InMux I__1199 (
            .O(N__5947),
            .I(N__5913));
    InMux I__1198 (
            .O(N__5946),
            .I(N__5913));
    InMux I__1197 (
            .O(N__5945),
            .I(N__5913));
    InMux I__1196 (
            .O(N__5944),
            .I(N__5908));
    InMux I__1195 (
            .O(N__5943),
            .I(N__5908));
    InMux I__1194 (
            .O(N__5942),
            .I(N__5903));
    InMux I__1193 (
            .O(N__5941),
            .I(N__5903));
    LocalMux I__1192 (
            .O(N__5936),
            .I(N__5865));
    InMux I__1191 (
            .O(N__5935),
            .I(N__5848));
    InMux I__1190 (
            .O(N__5934),
            .I(N__5848));
    InMux I__1189 (
            .O(N__5933),
            .I(N__5848));
    InMux I__1188 (
            .O(N__5932),
            .I(N__5848));
    InMux I__1187 (
            .O(N__5931),
            .I(N__5848));
    InMux I__1186 (
            .O(N__5930),
            .I(N__5848));
    InMux I__1185 (
            .O(N__5929),
            .I(N__5848));
    InMux I__1184 (
            .O(N__5928),
            .I(N__5848));
    InMux I__1183 (
            .O(N__5927),
            .I(N__5841));
    InMux I__1182 (
            .O(N__5926),
            .I(N__5841));
    InMux I__1181 (
            .O(N__5925),
            .I(N__5841));
    LocalMux I__1180 (
            .O(N__5922),
            .I(N__5826));
    LocalMux I__1179 (
            .O(N__5913),
            .I(N__5826));
    LocalMux I__1178 (
            .O(N__5908),
            .I(N__5826));
    LocalMux I__1177 (
            .O(N__5903),
            .I(N__5823));
    InMux I__1176 (
            .O(N__5902),
            .I(N__5808));
    InMux I__1175 (
            .O(N__5901),
            .I(N__5808));
    InMux I__1174 (
            .O(N__5900),
            .I(N__5808));
    InMux I__1173 (
            .O(N__5899),
            .I(N__5808));
    InMux I__1172 (
            .O(N__5898),
            .I(N__5808));
    InMux I__1171 (
            .O(N__5897),
            .I(N__5808));
    InMux I__1170 (
            .O(N__5896),
            .I(N__5808));
    InMux I__1169 (
            .O(N__5895),
            .I(N__5791));
    InMux I__1168 (
            .O(N__5894),
            .I(N__5791));
    InMux I__1167 (
            .O(N__5893),
            .I(N__5791));
    InMux I__1166 (
            .O(N__5892),
            .I(N__5791));
    InMux I__1165 (
            .O(N__5891),
            .I(N__5791));
    InMux I__1164 (
            .O(N__5890),
            .I(N__5791));
    InMux I__1163 (
            .O(N__5889),
            .I(N__5791));
    InMux I__1162 (
            .O(N__5888),
            .I(N__5791));
    InMux I__1161 (
            .O(N__5887),
            .I(N__5774));
    InMux I__1160 (
            .O(N__5886),
            .I(N__5774));
    InMux I__1159 (
            .O(N__5885),
            .I(N__5774));
    InMux I__1158 (
            .O(N__5884),
            .I(N__5774));
    InMux I__1157 (
            .O(N__5883),
            .I(N__5774));
    InMux I__1156 (
            .O(N__5882),
            .I(N__5774));
    InMux I__1155 (
            .O(N__5881),
            .I(N__5774));
    InMux I__1154 (
            .O(N__5880),
            .I(N__5774));
    InMux I__1153 (
            .O(N__5879),
            .I(N__5759));
    InMux I__1152 (
            .O(N__5878),
            .I(N__5759));
    InMux I__1151 (
            .O(N__5877),
            .I(N__5759));
    InMux I__1150 (
            .O(N__5876),
            .I(N__5759));
    InMux I__1149 (
            .O(N__5875),
            .I(N__5759));
    InMux I__1148 (
            .O(N__5874),
            .I(N__5759));
    InMux I__1147 (
            .O(N__5873),
            .I(N__5759));
    InMux I__1146 (
            .O(N__5872),
            .I(N__5750));
    InMux I__1145 (
            .O(N__5871),
            .I(N__5750));
    InMux I__1144 (
            .O(N__5870),
            .I(N__5750));
    InMux I__1143 (
            .O(N__5869),
            .I(N__5750));
    InMux I__1142 (
            .O(N__5868),
            .I(N__5747));
    Span4Mux_v I__1141 (
            .O(N__5865),
            .I(N__5740));
    LocalMux I__1140 (
            .O(N__5848),
            .I(N__5740));
    LocalMux I__1139 (
            .O(N__5841),
            .I(N__5740));
    InMux I__1138 (
            .O(N__5840),
            .I(N__5723));
    InMux I__1137 (
            .O(N__5839),
            .I(N__5723));
    InMux I__1136 (
            .O(N__5838),
            .I(N__5723));
    InMux I__1135 (
            .O(N__5837),
            .I(N__5723));
    InMux I__1134 (
            .O(N__5836),
            .I(N__5723));
    InMux I__1133 (
            .O(N__5835),
            .I(N__5723));
    InMux I__1132 (
            .O(N__5834),
            .I(N__5723));
    InMux I__1131 (
            .O(N__5833),
            .I(N__5723));
    Odrv4 I__1130 (
            .O(N__5826),
            .I(\DFT.aZ0Z_0 ));
    Odrv4 I__1129 (
            .O(N__5823),
            .I(\DFT.aZ0Z_0 ));
    LocalMux I__1128 (
            .O(N__5808),
            .I(\DFT.aZ0Z_0 ));
    LocalMux I__1127 (
            .O(N__5791),
            .I(\DFT.aZ0Z_0 ));
    LocalMux I__1126 (
            .O(N__5774),
            .I(\DFT.aZ0Z_0 ));
    LocalMux I__1125 (
            .O(N__5759),
            .I(\DFT.aZ0Z_0 ));
    LocalMux I__1124 (
            .O(N__5750),
            .I(\DFT.aZ0Z_0 ));
    LocalMux I__1123 (
            .O(N__5747),
            .I(\DFT.aZ0Z_0 ));
    Odrv4 I__1122 (
            .O(N__5740),
            .I(\DFT.aZ0Z_0 ));
    LocalMux I__1121 (
            .O(N__5723),
            .I(\DFT.aZ0Z_0 ));
    CascadeMux I__1120 (
            .O(N__5702),
            .I(N__5699));
    InMux I__1119 (
            .O(N__5699),
            .I(N__5696));
    LocalMux I__1118 (
            .O(N__5696),
            .I(N__5693));
    Span4Mux_h I__1117 (
            .O(N__5693),
            .I(N__5690));
    Odrv4 I__1116 (
            .O(N__5690),
            .I(\DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_0 ));
    InMux I__1115 (
            .O(N__5687),
            .I(N__5683));
    InMux I__1114 (
            .O(N__5686),
            .I(N__5680));
    LocalMux I__1113 (
            .O(N__5683),
            .I(N__5677));
    LocalMux I__1112 (
            .O(N__5680),
            .I(N__5674));
    Span4Mux_h I__1111 (
            .O(N__5677),
            .I(N__5671));
    Span4Mux_v I__1110 (
            .O(N__5674),
            .I(N__5668));
    Odrv4 I__1109 (
            .O(N__5671),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_CO ));
    Odrv4 I__1108 (
            .O(N__5668),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_CO ));
    InMux I__1107 (
            .O(N__5663),
            .I(N__5659));
    CascadeMux I__1106 (
            .O(N__5662),
            .I(N__5656));
    LocalMux I__1105 (
            .O(N__5659),
            .I(N__5653));
    InMux I__1104 (
            .O(N__5656),
            .I(N__5650));
    Span4Mux_h I__1103 (
            .O(N__5653),
            .I(N__5647));
    LocalMux I__1102 (
            .O(N__5650),
            .I(N__5644));
    Odrv4 I__1101 (
            .O(N__5647),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_823 ));
    Odrv4 I__1100 (
            .O(N__5644),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_823 ));
    CEMux I__1099 (
            .O(N__5639),
            .I(N__5635));
    CEMux I__1098 (
            .O(N__5638),
            .I(N__5629));
    LocalMux I__1097 (
            .O(N__5635),
            .I(N__5626));
    CEMux I__1096 (
            .O(N__5634),
            .I(N__5623));
    CEMux I__1095 (
            .O(N__5633),
            .I(N__5619));
    CEMux I__1094 (
            .O(N__5632),
            .I(N__5616));
    LocalMux I__1093 (
            .O(N__5629),
            .I(N__5609));
    Span4Mux_h I__1092 (
            .O(N__5626),
            .I(N__5609));
    LocalMux I__1091 (
            .O(N__5623),
            .I(N__5609));
    CEMux I__1090 (
            .O(N__5622),
            .I(N__5606));
    LocalMux I__1089 (
            .O(N__5619),
            .I(N__5601));
    LocalMux I__1088 (
            .O(N__5616),
            .I(N__5601));
    Span4Mux_v I__1087 (
            .O(N__5609),
            .I(N__5596));
    LocalMux I__1086 (
            .O(N__5606),
            .I(N__5596));
    Span4Mux_v I__1085 (
            .O(N__5601),
            .I(N__5593));
    Span4Mux_h I__1084 (
            .O(N__5596),
            .I(N__5590));
    Span4Mux_h I__1083 (
            .O(N__5593),
            .I(N__5587));
    Odrv4 I__1082 (
            .O(N__5590),
            .I(\DFT.un1_state_4_0 ));
    Odrv4 I__1081 (
            .O(N__5587),
            .I(\DFT.un1_state_4_0 ));
    InMux I__1080 (
            .O(N__5582),
            .I(N__5579));
    LocalMux I__1079 (
            .O(N__5579),
            .I(N__5576));
    Span4Mux_v I__1078 (
            .O(N__5576),
            .I(N__5573));
    Odrv4 I__1077 (
            .O(N__5573),
            .I(X_0__13));
    IoInMux I__1076 (
            .O(N__5570),
            .I(N__5567));
    LocalMux I__1075 (
            .O(N__5567),
            .I(N__5564));
    Span4Mux_s2_v I__1074 (
            .O(N__5564),
            .I(N__5561));
    Span4Mux_v I__1073 (
            .O(N__5561),
            .I(N__5558));
    Sp12to4 I__1072 (
            .O(N__5558),
            .I(N__5555));
    Span12Mux_s9_h I__1071 (
            .O(N__5555),
            .I(N__5552));
    Odrv12 I__1070 (
            .O(N__5552),
            .I(o_X_c_7));
    CascadeMux I__1069 (
            .O(N__5549),
            .I(N__5546));
    InMux I__1068 (
            .O(N__5546),
            .I(N__5543));
    LocalMux I__1067 (
            .O(N__5543),
            .I(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_0 ));
    CascadeMux I__1066 (
            .O(N__5540),
            .I(N__5537));
    InMux I__1065 (
            .O(N__5537),
            .I(N__5534));
    LocalMux I__1064 (
            .O(N__5534),
            .I(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_0 ));
    InMux I__1063 (
            .O(N__5531),
            .I(N__5528));
    LocalMux I__1062 (
            .O(N__5528),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_727_THRU_CO ));
    InMux I__1061 (
            .O(N__5525),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_727 ));
    InMux I__1060 (
            .O(N__5522),
            .I(N__5519));
    LocalMux I__1059 (
            .O(N__5519),
            .I(N__5516));
    Span4Mux_v I__1058 (
            .O(N__5516),
            .I(N__5513));
    Odrv4 I__1057 (
            .O(N__5513),
            .I(\DFT.multiplier.regsA_un3_result_cry_12_0_c_RNO ));
    InMux I__1056 (
            .O(N__5510),
            .I(N__5507));
    LocalMux I__1055 (
            .O(N__5507),
            .I(N__5504));
    Span4Mux_h I__1054 (
            .O(N__5504),
            .I(N__5501));
    Odrv4 I__1053 (
            .O(N__5501),
            .I(\DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_0 ));
    InMux I__1052 (
            .O(N__5498),
            .I(N__5495));
    LocalMux I__1051 (
            .O(N__5495),
            .I(N__5492));
    Odrv4 I__1050 (
            .O(N__5492),
            .I(\DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_2 ));
    InMux I__1049 (
            .O(N__5489),
            .I(N__5486));
    LocalMux I__1048 (
            .O(N__5486),
            .I(N__5483));
    Span4Mux_h I__1047 (
            .O(N__5483),
            .I(N__5480));
    Span4Mux_v I__1046 (
            .O(N__5480),
            .I(N__5477));
    Odrv4 I__1045 (
            .O(N__5477),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_897 ));
    InMux I__1044 (
            .O(N__5474),
            .I(N__5471));
    LocalMux I__1043 (
            .O(N__5471),
            .I(N__5468));
    Span4Mux_h I__1042 (
            .O(N__5468),
            .I(N__5465));
    Span4Mux_v I__1041 (
            .O(N__5465),
            .I(N__5462));
    Odrv4 I__1040 (
            .O(N__5462),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_898 ));
    InMux I__1039 (
            .O(N__5459),
            .I(\DFT.multiplier.regsA_un3_result_cry_2_2 ));
    CascadeMux I__1038 (
            .O(N__5456),
            .I(N__5453));
    InMux I__1037 (
            .O(N__5453),
            .I(N__5450));
    LocalMux I__1036 (
            .O(N__5450),
            .I(N__5447));
    Span4Mux_h I__1035 (
            .O(N__5447),
            .I(N__5444));
    Span4Mux_v I__1034 (
            .O(N__5444),
            .I(N__5441));
    Odrv4 I__1033 (
            .O(N__5441),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_899 ));
    InMux I__1032 (
            .O(N__5438),
            .I(\DFT.multiplier.regsA_un3_result_cry_3_1 ));
    CascadeMux I__1031 (
            .O(N__5435),
            .I(N__5432));
    InMux I__1030 (
            .O(N__5432),
            .I(N__5429));
    LocalMux I__1029 (
            .O(N__5429),
            .I(\DFT.multiplier.regsA_un3_result_6_a ));
    InMux I__1028 (
            .O(N__5426),
            .I(\DFT.multiplier.regsA_un3_result_cry_4 ));
    InMux I__1027 (
            .O(N__5423),
            .I(N__5420));
    LocalMux I__1026 (
            .O(N__5420),
            .I(N__5417));
    Odrv4 I__1025 (
            .O(N__5417),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_900 ));
    CascadeMux I__1024 (
            .O(N__5414),
            .I(N__5411));
    InMux I__1023 (
            .O(N__5411),
            .I(N__5408));
    LocalMux I__1022 (
            .O(N__5408),
            .I(N__5405));
    Odrv4 I__1021 (
            .O(N__5405),
            .I(\DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_0 ));
    InMux I__1020 (
            .O(N__5402),
            .I(N__5399));
    LocalMux I__1019 (
            .O(N__5399),
            .I(N__5396));
    Odrv4 I__1018 (
            .O(N__5396),
            .I(\DFT.multiplier.regsA_un3_result_5_b_l_ofx_1 ));
    CascadeMux I__1017 (
            .O(N__5393),
            .I(N__5390));
    InMux I__1016 (
            .O(N__5390),
            .I(N__5387));
    LocalMux I__1015 (
            .O(N__5387),
            .I(N__5384));
    Odrv4 I__1014 (
            .O(N__5384),
            .I(\DFT.multiplier.regsA_un3_result_cry_6_ma_0 ));
    InMux I__1013 (
            .O(N__5381),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_764 ));
    InMux I__1012 (
            .O(N__5378),
            .I(N__5375));
    LocalMux I__1011 (
            .O(N__5375),
            .I(N__5372));
    Span4Mux_h I__1010 (
            .O(N__5372),
            .I(N__5369));
    Odrv4 I__1009 (
            .O(N__5369),
            .I(\DFT.multiplier.regsA_un3_result_axb_3 ));
    InMux I__1008 (
            .O(N__5366),
            .I(N__5363));
    LocalMux I__1007 (
            .O(N__5363),
            .I(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO ));
    CascadeMux I__1006 (
            .O(N__5360),
            .I(N__5357));
    InMux I__1005 (
            .O(N__5357),
            .I(N__5354));
    LocalMux I__1004 (
            .O(N__5354),
            .I(N__5351));
    Odrv4 I__1003 (
            .O(N__5351),
            .I(\DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO_0 ));
    InMux I__1002 (
            .O(N__5348),
            .I(N__5345));
    LocalMux I__1001 (
            .O(N__5345),
            .I(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO ));
    InMux I__1000 (
            .O(N__5342),
            .I(N__5338));
    CascadeMux I__999 (
            .O(N__5341),
            .I(N__5335));
    LocalMux I__998 (
            .O(N__5338),
            .I(N__5332));
    InMux I__997 (
            .O(N__5335),
            .I(N__5329));
    Odrv4 I__996 (
            .O(N__5332),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_963 ));
    LocalMux I__995 (
            .O(N__5329),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_963 ));
    InMux I__994 (
            .O(N__5324),
            .I(N__5320));
    InMux I__993 (
            .O(N__5323),
            .I(N__5317));
    LocalMux I__992 (
            .O(N__5320),
            .I(\DFT.x_14 ));
    LocalMux I__991 (
            .O(N__5317),
            .I(\DFT.x_14 ));
    CascadeMux I__990 (
            .O(N__5312),
            .I(N__5309));
    InMux I__989 (
            .O(N__5309),
            .I(N__5305));
    InMux I__988 (
            .O(N__5308),
            .I(N__5302));
    LocalMux I__987 (
            .O(N__5305),
            .I(\DFT.x_11 ));
    LocalMux I__986 (
            .O(N__5302),
            .I(\DFT.x_11 ));
    InMux I__985 (
            .O(N__5297),
            .I(N__5294));
    LocalMux I__984 (
            .O(N__5294),
            .I(\DFT.multiplier.regsA_un3_result_cry_6_ma_2 ));
    CascadeMux I__983 (
            .O(N__5291),
            .I(N__5288));
    InMux I__982 (
            .O(N__5288),
            .I(N__5285));
    LocalMux I__981 (
            .O(N__5285),
            .I(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_5 ));
    CascadeMux I__980 (
            .O(N__5282),
            .I(N__5279));
    InMux I__979 (
            .O(N__5279),
            .I(N__5276));
    LocalMux I__978 (
            .O(N__5276),
            .I(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_4 ));
    CascadeMux I__977 (
            .O(N__5273),
            .I(N__5270));
    InMux I__976 (
            .O(N__5270),
            .I(N__5267));
    LocalMux I__975 (
            .O(N__5267),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_ma_3 ));
    CascadeMux I__974 (
            .O(N__5264),
            .I(N__5261));
    InMux I__973 (
            .O(N__5261),
            .I(N__5258));
    LocalMux I__972 (
            .O(N__5258),
            .I(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_4 ));
    CascadeMux I__971 (
            .O(N__5255),
            .I(N__5252));
    InMux I__970 (
            .O(N__5252),
            .I(N__5249));
    LocalMux I__969 (
            .O(N__5249),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_3 ));
    CascadeMux I__968 (
            .O(N__5246),
            .I(N__5243));
    InMux I__967 (
            .O(N__5243),
            .I(N__5240));
    LocalMux I__966 (
            .O(N__5240),
            .I(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_5 ));
    InMux I__965 (
            .O(N__5237),
            .I(N__5234));
    LocalMux I__964 (
            .O(N__5234),
            .I(N__5231));
    Span4Mux_h I__963 (
            .O(N__5231),
            .I(N__5228));
    Odrv4 I__962 (
            .O(N__5228),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_763_THRU_CO ));
    InMux I__961 (
            .O(N__5225),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_763 ));
    InMux I__960 (
            .O(N__5222),
            .I(N__5218));
    InMux I__959 (
            .O(N__5221),
            .I(N__5214));
    LocalMux I__958 (
            .O(N__5218),
            .I(N__5211));
    InMux I__957 (
            .O(N__5217),
            .I(N__5208));
    LocalMux I__956 (
            .O(N__5214),
            .I(N__5204));
    Span4Mux_h I__955 (
            .O(N__5211),
            .I(N__5201));
    LocalMux I__954 (
            .O(N__5208),
            .I(N__5198));
    InMux I__953 (
            .O(N__5207),
            .I(N__5195));
    Odrv4 I__952 (
            .O(N__5204),
            .I(\DFT.stateZ0Z_0 ));
    Odrv4 I__951 (
            .O(N__5201),
            .I(\DFT.stateZ0Z_0 ));
    Odrv12 I__950 (
            .O(N__5198),
            .I(\DFT.stateZ0Z_0 ));
    LocalMux I__949 (
            .O(N__5195),
            .I(\DFT.stateZ0Z_0 ));
    InMux I__948 (
            .O(N__5186),
            .I(N__5183));
    LocalMux I__947 (
            .O(N__5183),
            .I(N__5180));
    Span4Mux_v I__946 (
            .O(N__5180),
            .I(N__5175));
    InMux I__945 (
            .O(N__5179),
            .I(N__5172));
    InMux I__944 (
            .O(N__5178),
            .I(N__5168));
    Span4Mux_h I__943 (
            .O(N__5175),
            .I(N__5160));
    LocalMux I__942 (
            .O(N__5172),
            .I(N__5160));
    CascadeMux I__941 (
            .O(N__5171),
            .I(N__5157));
    LocalMux I__940 (
            .O(N__5168),
            .I(N__5154));
    InMux I__939 (
            .O(N__5167),
            .I(N__5147));
    InMux I__938 (
            .O(N__5166),
            .I(N__5147));
    InMux I__937 (
            .O(N__5165),
            .I(N__5147));
    Span4Mux_h I__936 (
            .O(N__5160),
            .I(N__5144));
    InMux I__935 (
            .O(N__5157),
            .I(N__5141));
    Span4Mux_v I__934 (
            .O(N__5154),
            .I(N__5138));
    LocalMux I__933 (
            .O(N__5147),
            .I(N__5135));
    Span4Mux_h I__932 (
            .O(N__5144),
            .I(N__5130));
    LocalMux I__931 (
            .O(N__5141),
            .I(N__5130));
    Span4Mux_h I__930 (
            .O(N__5138),
            .I(N__5125));
    Span4Mux_v I__929 (
            .O(N__5135),
            .I(N__5125));
    Span4Mux_v I__928 (
            .O(N__5130),
            .I(N__5122));
    Sp12to4 I__927 (
            .O(N__5125),
            .I(N__5119));
    Span4Mux_h I__926 (
            .O(N__5122),
            .I(N__5116));
    Span12Mux_h I__925 (
            .O(N__5119),
            .I(N__5111));
    Sp12to4 I__924 (
            .O(N__5116),
            .I(N__5111));
    Span12Mux_v I__923 (
            .O(N__5111),
            .I(N__5108));
    Odrv12 I__922 (
            .O(N__5108),
            .I(i_rst_c));
    CascadeMux I__921 (
            .O(N__5105),
            .I(N__5102));
    InMux I__920 (
            .O(N__5102),
            .I(N__5099));
    LocalMux I__919 (
            .O(N__5099),
            .I(\DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_1 ));
    InMux I__918 (
            .O(N__5096),
            .I(N__5093));
    LocalMux I__917 (
            .O(N__5093),
            .I(N__5088));
    InMux I__916 (
            .O(N__5092),
            .I(N__5083));
    InMux I__915 (
            .O(N__5091),
            .I(N__5083));
    Odrv4 I__914 (
            .O(N__5088),
            .I(\DFT.state_2_0 ));
    LocalMux I__913 (
            .O(N__5083),
            .I(\DFT.state_2_0 ));
    InMux I__912 (
            .O(N__5078),
            .I(N__5073));
    InMux I__911 (
            .O(N__5077),
            .I(N__5067));
    InMux I__910 (
            .O(N__5076),
            .I(N__5067));
    LocalMux I__909 (
            .O(N__5073),
            .I(N__5062));
    InMux I__908 (
            .O(N__5072),
            .I(N__5059));
    LocalMux I__907 (
            .O(N__5067),
            .I(N__5056));
    InMux I__906 (
            .O(N__5066),
            .I(N__5051));
    InMux I__905 (
            .O(N__5065),
            .I(N__5051));
    Span4Mux_h I__904 (
            .O(N__5062),
            .I(N__5048));
    LocalMux I__903 (
            .O(N__5059),
            .I(N__5045));
    Odrv4 I__902 (
            .O(N__5056),
            .I(\DFT.stateZ0Z_1 ));
    LocalMux I__901 (
            .O(N__5051),
            .I(\DFT.stateZ0Z_1 ));
    Odrv4 I__900 (
            .O(N__5048),
            .I(\DFT.stateZ0Z_1 ));
    Odrv12 I__899 (
            .O(N__5045),
            .I(\DFT.stateZ0Z_1 ));
    CascadeMux I__898 (
            .O(N__5036),
            .I(N__5033));
    InMux I__897 (
            .O(N__5033),
            .I(N__5030));
    LocalMux I__896 (
            .O(N__5030),
            .I(\DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_1 ));
    CascadeMux I__895 (
            .O(N__5027),
            .I(N__5024));
    InMux I__894 (
            .O(N__5024),
            .I(N__5021));
    LocalMux I__893 (
            .O(N__5021),
            .I(\DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_1 ));
    CascadeMux I__892 (
            .O(N__5018),
            .I(N__5015));
    InMux I__891 (
            .O(N__5015),
            .I(N__5012));
    LocalMux I__890 (
            .O(N__5012),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_ma_2 ));
    CascadeMux I__889 (
            .O(N__5009),
            .I(N__5006));
    InMux I__888 (
            .O(N__5006),
            .I(N__5003));
    LocalMux I__887 (
            .O(N__5003),
            .I(\DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO_0 ));
    InMux I__886 (
            .O(N__5000),
            .I(N__4997));
    LocalMux I__885 (
            .O(N__4997),
            .I(N__4994));
    Odrv4 I__884 (
            .O(N__4994),
            .I(\DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO ));
    InMux I__883 (
            .O(N__4991),
            .I(N__4988));
    LocalMux I__882 (
            .O(N__4988),
            .I(\DFT.multiplier.regsA_un3_result_5_b_l_ofx_2 ));
    InMux I__881 (
            .O(N__4985),
            .I(N__4982));
    LocalMux I__880 (
            .O(N__4982),
            .I(N__4979));
    Odrv4 I__879 (
            .O(N__4979),
            .I(X_0__15));
    IoInMux I__878 (
            .O(N__4976),
            .I(N__4972));
    IoInMux I__877 (
            .O(N__4975),
            .I(N__4969));
    LocalMux I__876 (
            .O(N__4972),
            .I(N__4963));
    LocalMux I__875 (
            .O(N__4969),
            .I(N__4963));
    IoInMux I__874 (
            .O(N__4968),
            .I(N__4960));
    IoSpan4Mux I__873 (
            .O(N__4963),
            .I(N__4955));
    LocalMux I__872 (
            .O(N__4960),
            .I(N__4952));
    IoInMux I__871 (
            .O(N__4959),
            .I(N__4949));
    IoInMux I__870 (
            .O(N__4958),
            .I(N__4946));
    IoSpan4Mux I__869 (
            .O(N__4955),
            .I(N__4939));
    IoSpan4Mux I__868 (
            .O(N__4952),
            .I(N__4939));
    LocalMux I__867 (
            .O(N__4949),
            .I(N__4939));
    LocalMux I__866 (
            .O(N__4946),
            .I(N__4934));
    IoSpan4Mux I__865 (
            .O(N__4939),
            .I(N__4931));
    IoInMux I__864 (
            .O(N__4938),
            .I(N__4928));
    IoInMux I__863 (
            .O(N__4937),
            .I(N__4925));
    IoSpan4Mux I__862 (
            .O(N__4934),
            .I(N__4922));
    Span4Mux_s3_v I__861 (
            .O(N__4931),
            .I(N__4919));
    LocalMux I__860 (
            .O(N__4928),
            .I(N__4916));
    LocalMux I__859 (
            .O(N__4925),
            .I(N__4913));
    IoSpan4Mux I__858 (
            .O(N__4922),
            .I(N__4910));
    Span4Mux_v I__857 (
            .O(N__4919),
            .I(N__4905));
    Span4Mux_s3_v I__856 (
            .O(N__4916),
            .I(N__4905));
    Span12Mux_s6_v I__855 (
            .O(N__4913),
            .I(N__4902));
    Span4Mux_s3_v I__854 (
            .O(N__4910),
            .I(N__4897));
    Span4Mux_h I__853 (
            .O(N__4905),
            .I(N__4897));
    Odrv12 I__852 (
            .O(N__4902),
            .I(o_X_c_15));
    Odrv4 I__851 (
            .O(N__4897),
            .I(o_X_c_15));
    CascadeMux I__850 (
            .O(N__4892),
            .I(N__4889));
    InMux I__849 (
            .O(N__4889),
            .I(N__4886));
    LocalMux I__848 (
            .O(N__4886),
            .I(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_3 ));
    CascadeMux I__847 (
            .O(N__4883),
            .I(N__4880));
    InMux I__846 (
            .O(N__4880),
            .I(N__4877));
    LocalMux I__845 (
            .O(N__4877),
            .I(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_3 ));
    CascadeMux I__844 (
            .O(N__4874),
            .I(N__4871));
    InMux I__843 (
            .O(N__4871),
            .I(N__4868));
    LocalMux I__842 (
            .O(N__4868),
            .I(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_4 ));
    CascadeMux I__841 (
            .O(N__4865),
            .I(N__4862));
    InMux I__840 (
            .O(N__4862),
            .I(N__4859));
    LocalMux I__839 (
            .O(N__4859),
            .I(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_4 ));
    CascadeMux I__838 (
            .O(N__4856),
            .I(N__4853));
    InMux I__837 (
            .O(N__4853),
            .I(N__4850));
    LocalMux I__836 (
            .O(N__4850),
            .I(N__4847));
    Odrv4 I__835 (
            .O(N__4847),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_1 ));
    CascadeMux I__834 (
            .O(N__4844),
            .I(N__4841));
    InMux I__833 (
            .O(N__4841),
            .I(N__4838));
    LocalMux I__832 (
            .O(N__4838),
            .I(\DFT.multiplier.regsA_un3_result_6_b_l_ofx ));
    InMux I__831 (
            .O(N__4835),
            .I(N__4832));
    LocalMux I__830 (
            .O(N__4832),
            .I(\DFT.multiplier.regsA_un3_result_cry_6_ma_1 ));
    CascadeMux I__829 (
            .O(N__4829),
            .I(N__4826));
    InMux I__828 (
            .O(N__4826),
            .I(N__4823));
    LocalMux I__827 (
            .O(N__4823),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_2 ));
    CascadeMux I__826 (
            .O(N__4820),
            .I(N__4817));
    InMux I__825 (
            .O(N__4817),
            .I(N__4814));
    LocalMux I__824 (
            .O(N__4814),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_965 ));
    InMux I__823 (
            .O(N__4811),
            .I(\DFT.multiplier.regsA_un3_result_cry_3 ));
    CascadeMux I__822 (
            .O(N__4808),
            .I(N__4805));
    InMux I__821 (
            .O(N__4805),
            .I(N__4802));
    LocalMux I__820 (
            .O(N__4802),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_966 ));
    InMux I__819 (
            .O(N__4799),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_0 ));
    InMux I__818 (
            .O(N__4796),
            .I(N__4793));
    LocalMux I__817 (
            .O(N__4793),
            .I(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNIRG904 ));
    CascadeMux I__816 (
            .O(N__4790),
            .I(N__4786));
    InMux I__815 (
            .O(N__4789),
            .I(N__4783));
    InMux I__814 (
            .O(N__4786),
            .I(N__4780));
    LocalMux I__813 (
            .O(N__4783),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_967 ));
    LocalMux I__812 (
            .O(N__4780),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_967 ));
    InMux I__811 (
            .O(N__4775),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_0 ));
    InMux I__810 (
            .O(N__4772),
            .I(N__4769));
    LocalMux I__809 (
            .O(N__4769),
            .I(\DFT.multiplier.regsA_un3_result_axb_7 ));
    InMux I__808 (
            .O(N__4766),
            .I(\DFT.multiplier.regsA_un3_result_cry_6_2 ));
    CEMux I__807 (
            .O(N__4763),
            .I(N__4759));
    CEMux I__806 (
            .O(N__4762),
            .I(N__4755));
    LocalMux I__805 (
            .O(N__4759),
            .I(N__4752));
    CEMux I__804 (
            .O(N__4758),
            .I(N__4747));
    LocalMux I__803 (
            .O(N__4755),
            .I(N__4744));
    Span4Mux_v I__802 (
            .O(N__4752),
            .I(N__4741));
    CEMux I__801 (
            .O(N__4751),
            .I(N__4738));
    CEMux I__800 (
            .O(N__4750),
            .I(N__4735));
    LocalMux I__799 (
            .O(N__4747),
            .I(N__4732));
    Span4Mux_v I__798 (
            .O(N__4744),
            .I(N__4725));
    Span4Mux_h I__797 (
            .O(N__4741),
            .I(N__4725));
    LocalMux I__796 (
            .O(N__4738),
            .I(N__4725));
    LocalMux I__795 (
            .O(N__4735),
            .I(N__4722));
    Span4Mux_h I__794 (
            .O(N__4732),
            .I(N__4719));
    Span4Mux_h I__793 (
            .O(N__4725),
            .I(N__4716));
    Span4Mux_h I__792 (
            .O(N__4722),
            .I(N__4713));
    Odrv4 I__791 (
            .O(N__4719),
            .I(\DFT.un1_state_1_0 ));
    Odrv4 I__790 (
            .O(N__4716),
            .I(\DFT.un1_state_1_0 ));
    Odrv4 I__789 (
            .O(N__4713),
            .I(\DFT.un1_state_1_0 ));
    InMux I__788 (
            .O(N__4706),
            .I(N__4702));
    InMux I__787 (
            .O(N__4705),
            .I(N__4699));
    LocalMux I__786 (
            .O(N__4702),
            .I(\DFT.x_13 ));
    LocalMux I__785 (
            .O(N__4699),
            .I(\DFT.x_13 ));
    InMux I__784 (
            .O(N__4694),
            .I(N__4690));
    InMux I__783 (
            .O(N__4693),
            .I(N__4687));
    LocalMux I__782 (
            .O(N__4690),
            .I(\DFT.x_12 ));
    LocalMux I__781 (
            .O(N__4687),
            .I(\DFT.x_12 ));
    InMux I__780 (
            .O(N__4682),
            .I(N__4678));
    InMux I__779 (
            .O(N__4681),
            .I(N__4675));
    LocalMux I__778 (
            .O(N__4678),
            .I(\DFT.x_15 ));
    LocalMux I__777 (
            .O(N__4675),
            .I(\DFT.x_15 ));
    InMux I__776 (
            .O(N__4670),
            .I(N__4667));
    LocalMux I__775 (
            .O(N__4667),
            .I(N__4664));
    Span4Mux_h I__774 (
            .O(N__4664),
            .I(N__4661));
    Odrv4 I__773 (
            .O(N__4661),
            .I(\DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO ));
    InMux I__772 (
            .O(N__4658),
            .I(N__4654));
    InMux I__771 (
            .O(N__4657),
            .I(N__4651));
    LocalMux I__770 (
            .O(N__4654),
            .I(\DFT.x_7 ));
    LocalMux I__769 (
            .O(N__4651),
            .I(\DFT.x_7 ));
    InMux I__768 (
            .O(N__4646),
            .I(N__4642));
    InMux I__767 (
            .O(N__4645),
            .I(N__4639));
    LocalMux I__766 (
            .O(N__4642),
            .I(\DFT.x_9 ));
    LocalMux I__765 (
            .O(N__4639),
            .I(\DFT.x_9 ));
    InMux I__764 (
            .O(N__4634),
            .I(N__4630));
    InMux I__763 (
            .O(N__4633),
            .I(N__4627));
    LocalMux I__762 (
            .O(N__4630),
            .I(\DFT.x_8 ));
    LocalMux I__761 (
            .O(N__4627),
            .I(\DFT.x_8 ));
    InMux I__760 (
            .O(N__4622),
            .I(\DFT.multiplier.regsA_un3_result_cry_2 ));
    CascadeMux I__759 (
            .O(N__4619),
            .I(N__4616));
    InMux I__758 (
            .O(N__4616),
            .I(N__4613));
    LocalMux I__757 (
            .O(N__4613),
            .I(N__4610));
    Span4Mux_h I__756 (
            .O(N__4610),
            .I(N__4607));
    Odrv4 I__755 (
            .O(N__4607),
            .I(\DFT.multiplier.regsA_un3_result_cry_2_THRU_CO ));
    InMux I__754 (
            .O(N__4604),
            .I(N__4601));
    LocalMux I__753 (
            .O(N__4601),
            .I(N__4598));
    Span4Mux_v I__752 (
            .O(N__4598),
            .I(N__4595));
    Odrv4 I__751 (
            .O(N__4595),
            .I(X_1__10));
    CascadeMux I__750 (
            .O(N__4592),
            .I(N__4589));
    InMux I__749 (
            .O(N__4589),
            .I(N__4586));
    LocalMux I__748 (
            .O(N__4586),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_964 ));
    InMux I__747 (
            .O(N__4583),
            .I(\DFT.multiplier.regsA_un3_result_cry_2_0 ));
    InMux I__746 (
            .O(N__4580),
            .I(N__4577));
    LocalMux I__745 (
            .O(N__4577),
            .I(N__4574));
    Odrv4 I__744 (
            .O(N__4574),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_659 ));
    InMux I__743 (
            .O(N__4571),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_7 ));
    CascadeMux I__742 (
            .O(N__4568),
            .I(N__4565));
    InMux I__741 (
            .O(N__4565),
            .I(N__4562));
    LocalMux I__740 (
            .O(N__4562),
            .I(N__4559));
    Odrv4 I__739 (
            .O(N__4559),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_660 ));
    InMux I__738 (
            .O(N__4556),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_7 ));
    InMux I__737 (
            .O(N__4553),
            .I(N__4550));
    LocalMux I__736 (
            .O(N__4550),
            .I(N__4547));
    Odrv4 I__735 (
            .O(N__4547),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_661_THRU_CO ));
    InMux I__734 (
            .O(N__4544),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_661 ));
    InMux I__733 (
            .O(N__4541),
            .I(bfn_11_20_0_));
    InMux I__732 (
            .O(N__4538),
            .I(N__4535));
    LocalMux I__731 (
            .O(N__4535),
            .I(N__4532));
    Odrv4 I__730 (
            .O(N__4532),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_662_THRU_CO ));
    InMux I__729 (
            .O(N__4529),
            .I(N__4526));
    LocalMux I__728 (
            .O(N__4526),
            .I(N__4523));
    Odrv4 I__727 (
            .O(N__4523),
            .I(\DFT.multiplier.regsA_un3_result_cry_13_0_c_RNO ));
    CascadeMux I__726 (
            .O(N__4520),
            .I(\DFT.state_2_0_cascade_ ));
    CascadeMux I__725 (
            .O(N__4517),
            .I(N__4514));
    InMux I__724 (
            .O(N__4514),
            .I(N__4511));
    LocalMux I__723 (
            .O(N__4511),
            .I(N__4508));
    Odrv4 I__722 (
            .O(N__4508),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_558_THRU_CO ));
    InMux I__721 (
            .O(N__4505),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_558 ));
    InMux I__720 (
            .O(N__4502),
            .I(N__4499));
    LocalMux I__719 (
            .O(N__4499),
            .I(N__4496));
    Odrv4 I__718 (
            .O(N__4496),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_559_THRU_CO ));
    InMux I__717 (
            .O(N__4493),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_559 ));
    InMux I__716 (
            .O(N__4490),
            .I(N__4487));
    LocalMux I__715 (
            .O(N__4487),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_594_THRU_CO ));
    InMux I__714 (
            .O(N__4484),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_560 ));
    InMux I__713 (
            .O(N__4481),
            .I(N__4478));
    LocalMux I__712 (
            .O(N__4478),
            .I(N__4475));
    Odrv4 I__711 (
            .O(N__4475),
            .I(\DFT.multiplier.regsA_un3_result_axb_13 ));
    CascadeMux I__710 (
            .O(N__4472),
            .I(N__4469));
    InMux I__709 (
            .O(N__4469),
            .I(N__4466));
    LocalMux I__708 (
            .O(N__4466),
            .I(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_3 ));
    InMux I__707 (
            .O(N__4463),
            .I(N__4457));
    InMux I__706 (
            .O(N__4462),
            .I(N__4457));
    LocalMux I__705 (
            .O(N__4457),
            .I(N__4454));
    Span4Mux_h I__704 (
            .O(N__4454),
            .I(N__4451));
    Odrv4 I__703 (
            .O(N__4451),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_655_THRU_CO ));
    InMux I__702 (
            .O(N__4448),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_655 ));
    InMux I__701 (
            .O(N__4445),
            .I(N__4442));
    LocalMux I__700 (
            .O(N__4442),
            .I(N__4439));
    Odrv4 I__699 (
            .O(N__4439),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_656_THRU_CO ));
    InMux I__698 (
            .O(N__4436),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_656 ));
    CascadeMux I__697 (
            .O(N__4433),
            .I(N__4430));
    InMux I__696 (
            .O(N__4430),
            .I(N__4427));
    LocalMux I__695 (
            .O(N__4427),
            .I(N__4424));
    Odrv4 I__694 (
            .O(N__4424),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_657_THRU_CO ));
    InMux I__693 (
            .O(N__4421),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_657 ));
    CascadeMux I__692 (
            .O(N__4418),
            .I(N__4415));
    InMux I__691 (
            .O(N__4415),
            .I(N__4412));
    LocalMux I__690 (
            .O(N__4412),
            .I(N__4409));
    Odrv4 I__689 (
            .O(N__4409),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_658_THRU_CO ));
    InMux I__688 (
            .O(N__4406),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_658 ));
    InMux I__687 (
            .O(N__4403),
            .I(N__4400));
    LocalMux I__686 (
            .O(N__4400),
            .I(N__4397));
    Span4Mux_h I__685 (
            .O(N__4397),
            .I(N__4394));
    Odrv4 I__684 (
            .O(N__4394),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_550_THRU_CO ));
    InMux I__683 (
            .O(N__4391),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_550 ));
    InMux I__682 (
            .O(N__4388),
            .I(N__4385));
    LocalMux I__681 (
            .O(N__4385),
            .I(N__4382));
    Odrv4 I__680 (
            .O(N__4382),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_551 ));
    InMux I__679 (
            .O(N__4379),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_6 ));
    InMux I__678 (
            .O(N__4376),
            .I(N__4373));
    LocalMux I__677 (
            .O(N__4373),
            .I(N__4370));
    Span4Mux_h I__676 (
            .O(N__4370),
            .I(N__4367));
    Odrv4 I__675 (
            .O(N__4367),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_552 ));
    InMux I__674 (
            .O(N__4364),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_6 ));
    InMux I__673 (
            .O(N__4361),
            .I(N__4358));
    LocalMux I__672 (
            .O(N__4358),
            .I(N__4355));
    Odrv4 I__671 (
            .O(N__4355),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_553_THRU_CO ));
    InMux I__670 (
            .O(N__4352),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_553 ));
    InMux I__669 (
            .O(N__4349),
            .I(N__4346));
    LocalMux I__668 (
            .O(N__4346),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_554_THRU_CO ));
    InMux I__667 (
            .O(N__4343),
            .I(bfn_11_18_0_));
    CascadeMux I__666 (
            .O(N__4340),
            .I(N__4337));
    InMux I__665 (
            .O(N__4337),
            .I(N__4334));
    LocalMux I__664 (
            .O(N__4334),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_555_THRU_CO ));
    InMux I__663 (
            .O(N__4331),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_555 ));
    InMux I__662 (
            .O(N__4328),
            .I(N__4325));
    LocalMux I__661 (
            .O(N__4325),
            .I(N__4322));
    Span4Mux_h I__660 (
            .O(N__4322),
            .I(N__4319));
    Odrv4 I__659 (
            .O(N__4319),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_556_THRU_CO ));
    InMux I__658 (
            .O(N__4316),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_556 ));
    InMux I__657 (
            .O(N__4313),
            .I(N__4310));
    LocalMux I__656 (
            .O(N__4310),
            .I(N__4307));
    Span4Mux_v I__655 (
            .O(N__4307),
            .I(N__4304));
    Odrv4 I__654 (
            .O(N__4304),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_557_THRU_CO ));
    InMux I__653 (
            .O(N__4301),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_557 ));
    InMux I__652 (
            .O(N__4298),
            .I(N__4295));
    LocalMux I__651 (
            .O(N__4295),
            .I(N__4292));
    Span4Mux_h I__650 (
            .O(N__4292),
            .I(N__4289));
    Odrv4 I__649 (
            .O(N__4289),
            .I(X_1__11));
    InMux I__648 (
            .O(N__4286),
            .I(N__4283));
    LocalMux I__647 (
            .O(N__4283),
            .I(X_1__13));
    InMux I__646 (
            .O(N__4280),
            .I(N__4277));
    LocalMux I__645 (
            .O(N__4277),
            .I(X_1__12));
    IoInMux I__644 (
            .O(N__4274),
            .I(N__4271));
    LocalMux I__643 (
            .O(N__4271),
            .I(N__4268));
    Span12Mux_s8_h I__642 (
            .O(N__4268),
            .I(N__4265));
    Odrv12 I__641 (
            .O(N__4265),
            .I(o_X_c_22));
    IoInMux I__640 (
            .O(N__4262),
            .I(N__4259));
    LocalMux I__639 (
            .O(N__4259),
            .I(N__4256));
    Span4Mux_s3_h I__638 (
            .O(N__4256),
            .I(N__4253));
    Span4Mux_h I__637 (
            .O(N__4253),
            .I(N__4250));
    Span4Mux_v I__636 (
            .O(N__4250),
            .I(N__4247));
    Odrv4 I__635 (
            .O(N__4247),
            .I(o_X_c_20));
    InMux I__634 (
            .O(N__4244),
            .I(N__4241));
    LocalMux I__633 (
            .O(N__4241),
            .I(N__4238));
    Span4Mux_v I__632 (
            .O(N__4238),
            .I(N__4235));
    Odrv4 I__631 (
            .O(N__4235),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_549_THRU_CO ));
    InMux I__630 (
            .O(N__4232),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_549 ));
    InMux I__629 (
            .O(N__4229),
            .I(N__4226));
    LocalMux I__628 (
            .O(N__4226),
            .I(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNI8J5C1 ));
    CascadeMux I__627 (
            .O(N__4223),
            .I(N__4219));
    InMux I__626 (
            .O(N__4222),
            .I(N__4216));
    InMux I__625 (
            .O(N__4219),
            .I(N__4213));
    LocalMux I__624 (
            .O(N__4216),
            .I(N__4208));
    LocalMux I__623 (
            .O(N__4213),
            .I(N__4208));
    Odrv4 I__622 (
            .O(N__4208),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_825 ));
    InMux I__621 (
            .O(N__4205),
            .I(\DFT.multiplier.regsA_un3_result_cry_3_0 ));
    InMux I__620 (
            .O(N__4202),
            .I(N__4199));
    LocalMux I__619 (
            .O(N__4199),
            .I(N__4196));
    Odrv4 I__618 (
            .O(N__4196),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_826 ));
    CascadeMux I__617 (
            .O(N__4193),
            .I(N__4190));
    InMux I__616 (
            .O(N__4190),
            .I(N__4187));
    LocalMux I__615 (
            .O(N__4187),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_860 ));
    InMux I__614 (
            .O(N__4184),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_8 ));
    InMux I__613 (
            .O(N__4181),
            .I(N__4178));
    LocalMux I__612 (
            .O(N__4178),
            .I(N__4175));
    Odrv12 I__611 (
            .O(N__4175),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_827 ));
    CascadeMux I__610 (
            .O(N__4172),
            .I(N__4169));
    InMux I__609 (
            .O(N__4169),
            .I(N__4166));
    LocalMux I__608 (
            .O(N__4166),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_861 ));
    InMux I__607 (
            .O(N__4163),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_1 ));
    InMux I__606 (
            .O(N__4160),
            .I(N__4157));
    LocalMux I__605 (
            .O(N__4157),
            .I(N__4154));
    Odrv4 I__604 (
            .O(N__4154),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_828 ));
    CascadeMux I__603 (
            .O(N__4151),
            .I(N__4148));
    InMux I__602 (
            .O(N__4148),
            .I(N__4145));
    LocalMux I__601 (
            .O(N__4145),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_862 ));
    InMux I__600 (
            .O(N__4142),
            .I(\DFT.multiplier.regsA_un3_result_cry_6 ));
    InMux I__599 (
            .O(N__4139),
            .I(N__4136));
    LocalMux I__598 (
            .O(N__4136),
            .I(N__4133));
    Odrv12 I__597 (
            .O(N__4133),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_829 ));
    CascadeMux I__596 (
            .O(N__4130),
            .I(N__4127));
    InMux I__595 (
            .O(N__4127),
            .I(N__4124));
    LocalMux I__594 (
            .O(N__4124),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_863 ));
    InMux I__593 (
            .O(N__4121),
            .I(\DFT.multiplier.regsA_un3_result_cry_7 ));
    InMux I__592 (
            .O(N__4118),
            .I(N__4115));
    LocalMux I__591 (
            .O(N__4115),
            .I(N__4112));
    Odrv12 I__590 (
            .O(N__4112),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_830 ));
    CascadeMux I__589 (
            .O(N__4109),
            .I(N__4106));
    InMux I__588 (
            .O(N__4106),
            .I(N__4103));
    LocalMux I__587 (
            .O(N__4103),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_864 ));
    InMux I__586 (
            .O(N__4100),
            .I(\DFT.multiplier.regsA_un3_result_cry_8_0 ));
    InMux I__585 (
            .O(N__4097),
            .I(N__4094));
    LocalMux I__584 (
            .O(N__4094),
            .I(N__4091));
    Odrv4 I__583 (
            .O(N__4091),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_831 ));
    CascadeMux I__582 (
            .O(N__4088),
            .I(N__4085));
    InMux I__581 (
            .O(N__4085),
            .I(N__4082));
    LocalMux I__580 (
            .O(N__4082),
            .I(N__4079));
    Odrv4 I__579 (
            .O(N__4079),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_865 ));
    InMux I__578 (
            .O(N__4076),
            .I(bfn_10_23_0_));
    InMux I__577 (
            .O(N__4073),
            .I(N__4070));
    LocalMux I__576 (
            .O(N__4070),
            .I(N__4067));
    Odrv4 I__575 (
            .O(N__4067),
            .I(\DFT.multiplier.regsA_un3_result_axb_11 ));
    InMux I__574 (
            .O(N__4064),
            .I(\DFT.multiplier.regsA_un3_result_cry_10 ));
    InMux I__573 (
            .O(N__4061),
            .I(N__4058));
    LocalMux I__572 (
            .O(N__4058),
            .I(N__4055));
    Odrv4 I__571 (
            .O(N__4055),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_623 ));
    InMux I__570 (
            .O(N__4052),
            .I(\DFT.multiplier.regsA_un3_result_cry_3_2 ));
    InMux I__569 (
            .O(N__4049),
            .I(N__4046));
    LocalMux I__568 (
            .O(N__4046),
            .I(N__4043));
    Odrv4 I__567 (
            .O(N__4043),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_624 ));
    InMux I__566 (
            .O(N__4040),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_1 ));
    CascadeMux I__565 (
            .O(N__4037),
            .I(N__4034));
    InMux I__564 (
            .O(N__4034),
            .I(N__4031));
    LocalMux I__563 (
            .O(N__4031),
            .I(N__4028));
    Odrv4 I__562 (
            .O(N__4028),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_625_THRU_CO ));
    InMux I__561 (
            .O(N__4025),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_2 ));
    InMux I__560 (
            .O(N__4022),
            .I(N__4019));
    LocalMux I__559 (
            .O(N__4019),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_626_THRU_CO ));
    InMux I__558 (
            .O(N__4016),
            .I(\DFT.multiplier.regsA_un3_result_cry_6_0 ));
    CascadeMux I__557 (
            .O(N__4013),
            .I(N__4010));
    InMux I__556 (
            .O(N__4010),
            .I(N__4007));
    LocalMux I__555 (
            .O(N__4007),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_627_THRU_CO ));
    InMux I__554 (
            .O(N__4004),
            .I(\DFT.multiplier.regsA_un3_result_cry_7_0 ));
    InMux I__553 (
            .O(N__4001),
            .I(\DFT.multiplier.regsA_un3_result_cry_8 ));
    InMux I__552 (
            .O(N__3998),
            .I(N__3995));
    LocalMux I__551 (
            .O(N__3995),
            .I(\DFT.multiplier.regsA_un3_result_cry_8_THRU_CO ));
    InMux I__550 (
            .O(N__3992),
            .I(N__3989));
    LocalMux I__549 (
            .O(N__3989),
            .I(N__3986));
    Odrv12 I__548 (
            .O(N__3986),
            .I(X_1__6));
    InMux I__547 (
            .O(N__3983),
            .I(N__3980));
    LocalMux I__546 (
            .O(N__3980),
            .I(N__3977));
    Span4Mux_h I__545 (
            .O(N__3977),
            .I(N__3974));
    Odrv4 I__544 (
            .O(N__3974),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_620_THRU_CO ));
    CascadeMux I__543 (
            .O(N__3971),
            .I(N__3968));
    InMux I__542 (
            .O(N__3968),
            .I(N__3965));
    LocalMux I__541 (
            .O(N__3965),
            .I(N__3962));
    Odrv12 I__540 (
            .O(N__3962),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_824 ));
    InMux I__539 (
            .O(N__3959),
            .I(\DFT.multiplier.regsA_un3_result_cry_2_1 ));
    CascadeMux I__538 (
            .O(N__3956),
            .I(N__3953));
    InMux I__537 (
            .O(N__3953),
            .I(N__3950));
    LocalMux I__536 (
            .O(N__3950),
            .I(N__3947));
    Odrv4 I__535 (
            .O(N__3947),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_588 ));
    InMux I__534 (
            .O(N__3944),
            .I(\DFT.multiplier.regsA_un3_result_cry_6_1 ));
    InMux I__533 (
            .O(N__3941),
            .I(N__3938));
    LocalMux I__532 (
            .O(N__3938),
            .I(N__3935));
    Odrv4 I__531 (
            .O(N__3935),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_589_THRU_CO ));
    InMux I__530 (
            .O(N__3932),
            .I(\DFT.multiplier.regsA_un3_result_cry_7_1 ));
    CascadeMux I__529 (
            .O(N__3929),
            .I(N__3926));
    InMux I__528 (
            .O(N__3926),
            .I(N__3923));
    LocalMux I__527 (
            .O(N__3923),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_590_THRU_CO ));
    InMux I__526 (
            .O(N__3920),
            .I(\DFT.multiplier.regsA_un3_result_cry_8_1 ));
    CascadeMux I__525 (
            .O(N__3917),
            .I(N__3914));
    InMux I__524 (
            .O(N__3914),
            .I(N__3911));
    LocalMux I__523 (
            .O(N__3911),
            .I(N__3908));
    Odrv4 I__522 (
            .O(N__3908),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_591_THRU_CO ));
    InMux I__521 (
            .O(N__3905),
            .I(bfn_10_20_0_));
    InMux I__520 (
            .O(N__3902),
            .I(N__3899));
    LocalMux I__519 (
            .O(N__3899),
            .I(N__3896));
    Odrv4 I__518 (
            .O(N__3896),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_592_THRU_CO ));
    InMux I__517 (
            .O(N__3893),
            .I(\DFT.multiplier.regsA_un3_result_cry_10_0 ));
    CascadeMux I__516 (
            .O(N__3890),
            .I(N__3887));
    InMux I__515 (
            .O(N__3887),
            .I(N__3884));
    LocalMux I__514 (
            .O(N__3884),
            .I(N__3881));
    Odrv4 I__513 (
            .O(N__3881),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_593_THRU_CO ));
    InMux I__512 (
            .O(N__3878),
            .I(\DFT.multiplier.regsA_un3_result_cry_11 ));
    CascadeMux I__511 (
            .O(N__3875),
            .I(N__3872));
    InMux I__510 (
            .O(N__3872),
            .I(N__3869));
    LocalMux I__509 (
            .O(N__3869),
            .I(\DFT.multiplier.regsA_un3_result_axb_9 ));
    InMux I__508 (
            .O(N__3866),
            .I(\DFT.multiplier.regsA_un3_result_cry_12 ));
    CascadeMux I__507 (
            .O(N__3863),
            .I(N__3860));
    InMux I__506 (
            .O(N__3860),
            .I(N__3857));
    LocalMux I__505 (
            .O(N__3857),
            .I(N__3854));
    Span4Mux_v I__504 (
            .O(N__3854),
            .I(N__3851));
    Odrv4 I__503 (
            .O(N__3851),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_621_THRU_CO ));
    CascadeMux I__502 (
            .O(N__3848),
            .I(N__3845));
    InMux I__501 (
            .O(N__3845),
            .I(N__3842));
    LocalMux I__500 (
            .O(N__3842),
            .I(N__3839));
    Odrv4 I__499 (
            .O(N__3839),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_622_THRU_CO ));
    InMux I__498 (
            .O(N__3836),
            .I(\DFT.multiplier.regsA_un3_result_cry_2_3 ));
    CascadeMux I__497 (
            .O(N__3833),
            .I(N__3830));
    InMux I__496 (
            .O(N__3830),
            .I(N__3827));
    LocalMux I__495 (
            .O(N__3827),
            .I(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_2 ));
    CascadeMux I__494 (
            .O(N__3824),
            .I(N__3821));
    InMux I__493 (
            .O(N__3821),
            .I(N__3818));
    LocalMux I__492 (
            .O(N__3818),
            .I(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_3 ));
    CascadeMux I__491 (
            .O(N__3815),
            .I(N__3812));
    InMux I__490 (
            .O(N__3812),
            .I(N__3809));
    LocalMux I__489 (
            .O(N__3809),
            .I(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_2 ));
    CascadeMux I__488 (
            .O(N__3806),
            .I(N__3803));
    InMux I__487 (
            .O(N__3803),
            .I(N__3800));
    LocalMux I__486 (
            .O(N__3800),
            .I(N__3797));
    Odrv4 I__485 (
            .O(N__3797),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_583_THRU_CO ));
    CascadeMux I__484 (
            .O(N__3794),
            .I(N__3791));
    InMux I__483 (
            .O(N__3791),
            .I(N__3788));
    LocalMux I__482 (
            .O(N__3788),
            .I(N__3785));
    Odrv4 I__481 (
            .O(N__3785),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_584_THRU_CO ));
    CascadeMux I__480 (
            .O(N__3782),
            .I(N__3779));
    InMux I__479 (
            .O(N__3779),
            .I(N__3776));
    LocalMux I__478 (
            .O(N__3776),
            .I(N__3773));
    Odrv4 I__477 (
            .O(N__3773),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_585_THRU_CO ));
    InMux I__476 (
            .O(N__3770),
            .I(\DFT.multiplier.regsA_un3_result_cry_3_3 ));
    CascadeMux I__475 (
            .O(N__3767),
            .I(N__3764));
    InMux I__474 (
            .O(N__3764),
            .I(N__3761));
    LocalMux I__473 (
            .O(N__3761),
            .I(N__3758));
    Odrv12 I__472 (
            .O(N__3758),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_586_THRU_CO ));
    InMux I__471 (
            .O(N__3755),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_2 ));
    CascadeMux I__470 (
            .O(N__3752),
            .I(N__3749));
    InMux I__469 (
            .O(N__3749),
            .I(N__3746));
    LocalMux I__468 (
            .O(N__3746),
            .I(N__3743));
    Odrv4 I__467 (
            .O(N__3743),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_587 ));
    InMux I__466 (
            .O(N__3740),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_3 ));
    InMux I__465 (
            .O(N__3737),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_586 ));
    CascadeMux I__464 (
            .O(N__3734),
            .I(N__3731));
    InMux I__463 (
            .O(N__3731),
            .I(N__3728));
    LocalMux I__462 (
            .O(N__3728),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_ma_1 ));
    InMux I__461 (
            .O(N__3725),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_5 ));
    InMux I__460 (
            .O(N__3722),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_5 ));
    InMux I__459 (
            .O(N__3719),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_589 ));
    InMux I__458 (
            .O(N__3716),
            .I(bfn_10_18_0_));
    InMux I__457 (
            .O(N__3713),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_591 ));
    InMux I__456 (
            .O(N__3710),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_592 ));
    InMux I__455 (
            .O(N__3707),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_593 ));
    InMux I__454 (
            .O(N__3704),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_594 ));
    InMux I__453 (
            .O(N__3701),
            .I(N__3698));
    LocalMux I__452 (
            .O(N__3698),
            .I(N__3695));
    Odrv4 I__451 (
            .O(N__3695),
            .I(X_1__8));
    InMux I__450 (
            .O(N__3692),
            .I(N__3689));
    LocalMux I__449 (
            .O(N__3689),
            .I(N__3686));
    Odrv4 I__448 (
            .O(N__3686),
            .I(X_1__9));
    InMux I__447 (
            .O(N__3683),
            .I(N__3680));
    LocalMux I__446 (
            .O(N__3680),
            .I(X_1__7));
    IoInMux I__445 (
            .O(N__3677),
            .I(N__3674));
    LocalMux I__444 (
            .O(N__3674),
            .I(N__3671));
    Span4Mux_s0_v I__443 (
            .O(N__3671),
            .I(N__3668));
    Sp12to4 I__442 (
            .O(N__3668),
            .I(N__3665));
    Span12Mux_s8_h I__441 (
            .O(N__3665),
            .I(N__3662));
    Odrv12 I__440 (
            .O(N__3662),
            .I(o_X_c_17));
    IoInMux I__439 (
            .O(N__3659),
            .I(N__3656));
    LocalMux I__438 (
            .O(N__3656),
            .I(N__3653));
    IoSpan4Mux I__437 (
            .O(N__3653),
            .I(N__3650));
    Span4Mux_s3_h I__436 (
            .O(N__3650),
            .I(N__3647));
    Span4Mux_h I__435 (
            .O(N__3647),
            .I(N__3644));
    Odrv4 I__434 (
            .O(N__3644),
            .I(o_X_c_23));
    InMux I__433 (
            .O(N__3641),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_583 ));
    InMux I__432 (
            .O(N__3638),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_584 ));
    InMux I__431 (
            .O(N__3635),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_585 ));
    CascadeMux I__430 (
            .O(N__3632),
            .I(N__3629));
    InMux I__429 (
            .O(N__3629),
            .I(N__3626));
    LocalMux I__428 (
            .O(N__3626),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_0 ));
    InMux I__427 (
            .O(N__3623),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_622 ));
    CascadeMux I__426 (
            .O(N__3620),
            .I(N__3617));
    InMux I__425 (
            .O(N__3617),
            .I(N__3614));
    LocalMux I__424 (
            .O(N__3614),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_ma_0 ));
    InMux I__423 (
            .O(N__3611),
            .I(\DFT.multiplier.regsA_un3_result_cry_4_4 ));
    InMux I__422 (
            .O(N__3608),
            .I(\DFT.multiplier.regsA_un3_result_cry_5_4 ));
    InMux I__421 (
            .O(N__3605),
            .I(N__3602));
    LocalMux I__420 (
            .O(N__3602),
            .I(\DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO ));
    InMux I__419 (
            .O(N__3599),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_625 ));
    InMux I__418 (
            .O(N__3596),
            .I(bfn_9_20_0_));
    InMux I__417 (
            .O(N__3593),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_627 ));
    InMux I__416 (
            .O(N__3590),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_628 ));
    InMux I__415 (
            .O(N__3587),
            .I(N__3584));
    LocalMux I__414 (
            .O(N__3584),
            .I(\DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO ));
    InMux I__413 (
            .O(N__3581),
            .I(N__3578));
    LocalMux I__412 (
            .O(N__3578),
            .I(\DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO ));
    CascadeMux I__411 (
            .O(N__3575),
            .I(N__3572));
    InMux I__410 (
            .O(N__3572),
            .I(N__3569));
    LocalMux I__409 (
            .O(N__3569),
            .I(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_2 ));
    CascadeMux I__408 (
            .O(N__3566),
            .I(N__3563));
    InMux I__407 (
            .O(N__3563),
            .I(N__3560));
    LocalMux I__406 (
            .O(N__3560),
            .I(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_2 ));
    InMux I__405 (
            .O(N__3557),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_619 ));
    CascadeMux I__404 (
            .O(N__3554),
            .I(N__3551));
    InMux I__403 (
            .O(N__3551),
            .I(N__3548));
    LocalMux I__402 (
            .O(N__3548),
            .I(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_1 ));
    InMux I__401 (
            .O(N__3545),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_620 ));
    CascadeMux I__400 (
            .O(N__3542),
            .I(N__3539));
    InMux I__399 (
            .O(N__3539),
            .I(N__3536));
    LocalMux I__398 (
            .O(N__3536),
            .I(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_1 ));
    InMux I__397 (
            .O(N__3533),
            .I(\DFT.multiplier.mult1_AdderTree2i_bigtree_621 ));
    CascadeMux I__396 (
            .O(N__3530),
            .I(\DFT.o_done_RNOZ0Z_0_cascade_ ));
    IoInMux I__395 (
            .O(N__3527),
            .I(N__3524));
    LocalMux I__394 (
            .O(N__3524),
            .I(N__3521));
    IoSpan4Mux I__393 (
            .O(N__3521),
            .I(N__3518));
    IoSpan4Mux I__392 (
            .O(N__3518),
            .I(N__3515));
    IoSpan4Mux I__391 (
            .O(N__3515),
            .I(N__3511));
    InMux I__390 (
            .O(N__3514),
            .I(N__3508));
    IoSpan4Mux I__389 (
            .O(N__3511),
            .I(N__3505));
    LocalMux I__388 (
            .O(N__3508),
            .I(N__3502));
    Span4Mux_s1_h I__387 (
            .O(N__3505),
            .I(N__3496));
    Span4Mux_v I__386 (
            .O(N__3502),
            .I(N__3496));
    InMux I__385 (
            .O(N__3501),
            .I(N__3493));
    Span4Mux_h I__384 (
            .O(N__3496),
            .I(N__3490));
    LocalMux I__383 (
            .O(N__3493),
            .I(done_c));
    Odrv4 I__382 (
            .O(N__3490),
            .I(done_c));
    InMux I__381 (
            .O(N__3485),
            .I(N__3482));
    LocalMux I__380 (
            .O(N__3482),
            .I(N__3478));
    InMux I__379 (
            .O(N__3481),
            .I(N__3475));
    Odrv4 I__378 (
            .O(N__3478),
            .I(\DFT.state_RNIHM3GZ0Z_0 ));
    LocalMux I__377 (
            .O(N__3475),
            .I(\DFT.state_RNIHM3GZ0Z_0 ));
    IoInMux I__376 (
            .O(N__3470),
            .I(N__3467));
    LocalMux I__375 (
            .O(N__3467),
            .I(N__3464));
    IoSpan4Mux I__374 (
            .O(N__3464),
            .I(N__3461));
    Span4Mux_s2_h I__373 (
            .O(N__3461),
            .I(N__3458));
    Span4Mux_h I__372 (
            .O(N__3458),
            .I(N__3455));
    Odrv4 I__371 (
            .O(N__3455),
            .I(o_X_c_18));
    IoInMux I__370 (
            .O(N__3452),
            .I(N__3449));
    LocalMux I__369 (
            .O(N__3449),
            .I(N__3446));
    IoSpan4Mux I__368 (
            .O(N__3446),
            .I(N__3443));
    Span4Mux_s3_v I__367 (
            .O(N__3443),
            .I(N__3440));
    Span4Mux_v I__366 (
            .O(N__3440),
            .I(N__3437));
    Odrv4 I__365 (
            .O(N__3437),
            .I(o_X_c_16));
    IoInMux I__364 (
            .O(N__3434),
            .I(N__3431));
    LocalMux I__363 (
            .O(N__3431),
            .I(N__3428));
    Span4Mux_s3_h I__362 (
            .O(N__3428),
            .I(N__3425));
    Span4Mux_v I__361 (
            .O(N__3425),
            .I(N__3422));
    Odrv4 I__360 (
            .O(N__3422),
            .I(o_X_c_19));
    IoInMux I__359 (
            .O(N__3419),
            .I(N__3416));
    LocalMux I__358 (
            .O(N__3416),
            .I(N__3413));
    IoSpan4Mux I__357 (
            .O(N__3413),
            .I(N__3410));
    Span4Mux_s2_h I__356 (
            .O(N__3410),
            .I(N__3407));
    Span4Mux_h I__355 (
            .O(N__3407),
            .I(N__3404));
    Odrv4 I__354 (
            .O(N__3404),
            .I(o_X_c_21));
    IoInMux I__353 (
            .O(N__3401),
            .I(N__3398));
    LocalMux I__352 (
            .O(N__3398),
            .I(N__3395));
    IoSpan4Mux I__351 (
            .O(N__3395),
            .I(N__3392));
    Span4Mux_s1_v I__350 (
            .O(N__3392),
            .I(N__3389));
    Sp12to4 I__349 (
            .O(N__3389),
            .I(N__3386));
    Span12Mux_s9_v I__348 (
            .O(N__3386),
            .I(N__3383));
    Span12Mux_v I__347 (
            .O(N__3383),
            .I(N__3380));
    Odrv12 I__346 (
            .O(N__3380),
            .I(i_ref_clk_c));
    IoInMux I__345 (
            .O(N__3377),
            .I(N__3374));
    LocalMux I__344 (
            .O(N__3374),
            .I(i_rst_c_i));
    IoInMux I__343 (
            .O(N__3371),
            .I(N__3368));
    LocalMux I__342 (
            .O(N__3368),
            .I(\DFT.done_c_0 ));
    ClkMux I__341 (
            .O(N__3365),
            .I(N__3278));
    ClkMux I__340 (
            .O(N__3364),
            .I(N__3278));
    ClkMux I__339 (
            .O(N__3363),
            .I(N__3278));
    ClkMux I__338 (
            .O(N__3362),
            .I(N__3278));
    ClkMux I__337 (
            .O(N__3361),
            .I(N__3278));
    ClkMux I__336 (
            .O(N__3360),
            .I(N__3278));
    ClkMux I__335 (
            .O(N__3359),
            .I(N__3278));
    ClkMux I__334 (
            .O(N__3358),
            .I(N__3278));
    ClkMux I__333 (
            .O(N__3357),
            .I(N__3278));
    ClkMux I__332 (
            .O(N__3356),
            .I(N__3278));
    ClkMux I__331 (
            .O(N__3355),
            .I(N__3278));
    ClkMux I__330 (
            .O(N__3354),
            .I(N__3278));
    ClkMux I__329 (
            .O(N__3353),
            .I(N__3278));
    ClkMux I__328 (
            .O(N__3352),
            .I(N__3278));
    ClkMux I__327 (
            .O(N__3351),
            .I(N__3278));
    ClkMux I__326 (
            .O(N__3350),
            .I(N__3278));
    ClkMux I__325 (
            .O(N__3349),
            .I(N__3278));
    ClkMux I__324 (
            .O(N__3348),
            .I(N__3278));
    ClkMux I__323 (
            .O(N__3347),
            .I(N__3278));
    ClkMux I__322 (
            .O(N__3346),
            .I(N__3278));
    ClkMux I__321 (
            .O(N__3345),
            .I(N__3278));
    ClkMux I__320 (
            .O(N__3344),
            .I(N__3278));
    ClkMux I__319 (
            .O(N__3343),
            .I(N__3278));
    ClkMux I__318 (
            .O(N__3342),
            .I(N__3278));
    ClkMux I__317 (
            .O(N__3341),
            .I(N__3278));
    ClkMux I__316 (
            .O(N__3340),
            .I(N__3278));
    ClkMux I__315 (
            .O(N__3339),
            .I(N__3278));
    ClkMux I__314 (
            .O(N__3338),
            .I(N__3278));
    ClkMux I__313 (
            .O(N__3337),
            .I(N__3278));
    GlobalMux I__312 (
            .O(N__3278),
            .I(N__3275));
    gio2CtrlBuf I__311 (
            .O(N__3275),
            .I(sys_clk_g));
    IoInMux I__310 (
            .O(N__3272),
            .I(N__3269));
    LocalMux I__309 (
            .O(N__3269),
            .I(N__3266));
    Odrv4 I__308 (
            .O(N__3266),
            .I(sys_clk));
    INV INVo_X_0__nesr_5C (
            .O(INVo_X_0__nesr_5C_net),
            .I(N__3338));
    INV INVo_X_1__nesr_9C (
            .O(INVo_X_1__nesr_9C_net),
            .I(N__3342));
    INV INVo_X_0__nesr_8C (
            .O(INVo_X_0__nesr_8C_net),
            .I(N__3339));
    INV INVo_X_0__nesr_4C (
            .O(INVo_X_0__nesr_4C_net),
            .I(N__3341));
    INV INVo_X_0__nesr_3C (
            .O(INVo_X_0__nesr_3C_net),
            .I(N__3348));
    INV INVo_X_1__nesr_8C (
            .O(INVo_X_1__nesr_8C_net),
            .I(N__3352));
    INV INVo_X_0__nesr_1C (
            .O(INVo_X_0__nesr_1C_net),
            .I(N__3354));
    INV INVo_X_0__nesr_7C (
            .O(INVo_X_0__nesr_7C_net),
            .I(N__3337));
    INV \INVDFT.o_X_0__nesr_6C  (
            .O(\INVDFT.o_X_0__nesr_6C_net ),
            .I(N__3353));
    INV \INVDFT.o_X_0__nesr_11C  (
            .O(\INVDFT.o_X_0__nesr_11C_net ),
            .I(N__3344));
    INV \INVDFT.o_X_0__nesr_14C  (
            .O(\INVDFT.o_X_0__nesr_14C_net ),
            .I(N__3347));
    INV \INVDFT.o_X_0__nesr_10C  (
            .O(\INVDFT.o_X_0__nesr_10C_net ),
            .I(N__3351));
    INV \INVDFT.b_6C  (
            .O(\INVDFT.b_6C_net ),
            .I(N__3362));
    INV INVo_X_0__nesr_9C (
            .O(INVo_X_0__nesr_9C_net),
            .I(N__3340));
    INV \INVDFT.o_X_0__nesr_13C  (
            .O(\INVDFT.o_X_0__nesr_13C_net ),
            .I(N__3346));
    INV \INVDFT.o_X_1__nesr_10C  (
            .O(\INVDFT.o_X_1__nesr_10C_net ),
            .I(N__3350));
    INV \INVDFT.o_X_0__nesr_7C  (
            .O(\INVDFT.o_X_0__nesr_7C_net ),
            .I(N__3357));
    INV \INVDFT.state_0C  (
            .O(\INVDFT.state_0C_net ),
            .I(N__3360));
    INV INVo_X_1__nesr_4C (
            .O(INVo_X_1__nesr_4C_net),
            .I(N__3343));
    INV INVo_X_1__nesr_6C (
            .O(INVo_X_1__nesr_6C_net),
            .I(N__3345));
    INV \INVDFT.o_X_1__nesr_12C  (
            .O(\INVDFT.o_X_1__nesr_12C_net ),
            .I(N__3349));
    INV \INVDFT.o_X_1__nesr_6C  (
            .O(\INVDFT.o_X_1__nesr_6C_net ),
            .I(N__3356));
    INV INVo_X_1__nesr_1C (
            .O(INVo_X_1__nesr_1C_net),
            .I(N__3355));
    INV \INVDFT.o_X_1__nesr_7C  (
            .O(\INVDFT.o_X_1__nesr_7C_net ),
            .I(N__3359));
    INV \INVDFT.o_X_1__nesr_8C  (
            .O(\INVDFT.o_X_1__nesr_8C_net ),
            .I(N__3361));
    INV INVo_X_1__nesr_5C (
            .O(INVo_X_1__nesr_5C_net),
            .I(N__3358));
    INV INVo_X_1__nesr_3C (
            .O(INVo_X_1__nesr_3C_net),
            .I(N__3363));
    INV INVo_X_1__nesr_2C (
            .O(INVo_X_1__nesr_2C_net),
            .I(N__3364));
    INV \INVDFT.o_doneC  (
            .O(\INVDFT.o_doneC_net ),
            .I(N__3365));
    defparam IN_MUX_bfv_10_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_19_0_));
    defparam IN_MUX_bfv_10_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_20_0_ (
            .carryinitin(\DFT.multiplier.regsA_un3_result_cry_9_0 ),
            .carryinitout(bfn_10_20_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_14_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_17_0_));
    defparam IN_MUX_bfv_14_18_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_14_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_14_18_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_11_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_20_0_ (
            .carryinitin(\DFT.multiplier.mult1_AdderTree2i_bigtree_662 ),
            .carryinitout(bfn_11_20_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_9_20_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_20_0_ (
            .carryinitin(\DFT.multiplier.mult1_AdderTree2i_bigtree_626 ),
            .carryinitout(bfn_9_20_0_));
    defparam IN_MUX_bfv_10_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_17_0_));
    defparam IN_MUX_bfv_10_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_18_0_ (
            .carryinitin(\DFT.multiplier.mult1_AdderTree2i_bigtree_590 ),
            .carryinitout(bfn_10_18_0_));
    defparam IN_MUX_bfv_11_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_17_0_));
    defparam IN_MUX_bfv_11_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_18_0_ (
            .carryinitin(\DFT.multiplier.mult1_AdderTree2i_bigtree_554 ),
            .carryinitout(bfn_11_18_0_));
    defparam IN_MUX_bfv_11_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_22_0_));
    defparam IN_MUX_bfv_13_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_17_0_));
    defparam IN_MUX_bfv_11_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_23_0_));
    defparam IN_MUX_bfv_10_21_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_21_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_21_0_));
    defparam IN_MUX_bfv_10_22_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_10_22_0_));
    defparam IN_MUX_bfv_10_23_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_10_23_0_ (
            .carryinitin(\DFT.multiplier.regsA_un3_result_cry_9 ),
            .carryinitout(bfn_10_23_0_));
    ICE_GB \DFT.o_done_RNI6TUH_0  (
            .USERSIGNALTOGLOBALBUFFER(N__3371),
            .GLOBALBUFFEROUTPUT(done_c_0_g));
    ICE_GB sys_clk_derived_clock_RNI5LTF (
            .USERSIGNALTOGLOBALBUFFER(N__3272),
            .GLOBALBUFFEROUTPUT(sys_clk_g));
    ICE_GB i_rst_ibuf_RNI6EKC_0 (
            .USERSIGNALTOGLOBALBUFFER(N__3377),
            .GLOBALBUFFEROUTPUT(i_rst_c_i_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam i_rst_ibuf_RNI6EKC_LC_1_16_3.C_ON=1'b0;
    defparam i_rst_ibuf_RNI6EKC_LC_1_16_3.SEQ_MODE=4'b0000;
    defparam i_rst_ibuf_RNI6EKC_LC_1_16_3.LUT_INIT=16'b0101010101010101;
    LogicCell40 i_rst_ibuf_RNI6EKC_LC_1_16_3 (
            .in0(N__5186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(i_rst_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.o_done_RNI6TUH_LC_1_17_2 .C_ON=1'b0;
    defparam \DFT.o_done_RNI6TUH_LC_1_17_2 .SEQ_MODE=4'b0000;
    defparam \DFT.o_done_RNI6TUH_LC_1_17_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \DFT.o_done_RNI6TUH_LC_1_17_2  (
            .in0(N__6528),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3514),
            .lcout(\DFT.done_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.o_done_RNO_0_LC_7_19_2 .C_ON=1'b0;
    defparam \DFT.o_done_RNO_0_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \DFT.o_done_RNO_0_LC_7_19_2 .LUT_INIT=16'b0101010101110111;
    LogicCell40 \DFT.o_done_RNO_0_LC_7_19_2  (
            .in0(N__5179),
            .in1(N__5222),
            .in2(_gnd_net_),
            .in3(N__5078),
            .lcout(),
            .ltout(\DFT.o_done_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.o_done_LC_7_19_3 .C_ON=1'b0;
    defparam \DFT.o_done_LC_7_19_3 .SEQ_MODE=4'b1000;
    defparam \DFT.o_done_LC_7_19_3 .LUT_INIT=16'b0000111100001100;
    LogicCell40 \DFT.o_done_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__3485),
            .in2(N__3530),
            .in3(N__3501),
            .lcout(done_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_doneC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.state_RNIHM3G_0_LC_7_20_3 .C_ON=1'b0;
    defparam \DFT.state_RNIHM3G_0_LC_7_20_3 .SEQ_MODE=4'b0000;
    defparam \DFT.state_RNIHM3G_0_LC_7_20_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \DFT.state_RNIHM3G_0_LC_7_20_3  (
            .in0(N__5178),
            .in1(N__5217),
            .in2(_gnd_net_),
            .in3(N__5072),
            .lcout(\DFT.state_RNIHM3GZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.state_RNIN4OS_0_LC_7_21_1 .C_ON=1'b0;
    defparam \DFT.state_RNIN4OS_0_LC_7_21_1 .SEQ_MODE=4'b0000;
    defparam \DFT.state_RNIN4OS_0_LC_7_21_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DFT.state_RNIN4OS_0_LC_7_21_1  (
            .in0(_gnd_net_),
            .in1(N__6529),
            .in2(_gnd_net_),
            .in3(N__3481),
            .lcout(\DFT.un1_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_X_1__nesr_2_LC_7_22_1.C_ON=1'b0;
    defparam o_X_1__nesr_2_LC_7_22_1.SEQ_MODE=4'b1000;
    defparam o_X_1__nesr_2_LC_7_22_1.LUT_INIT=16'b1100110011001100;
    LogicCell40 o_X_1__nesr_2_LC_7_22_1 (
            .in0(_gnd_net_),
            .in1(N__3701),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(o_X_c_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_1__nesr_2C_net),
            .ce(N__6567),
            .sr(N__6490));
    defparam o_X_1__nesr_0_LC_7_22_3.C_ON=1'b0;
    defparam o_X_1__nesr_0_LC_7_22_3.SEQ_MODE=4'b1000;
    defparam o_X_1__nesr_0_LC_7_22_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_1__nesr_0_LC_7_22_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3992),
            .lcout(o_X_c_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_1__nesr_2C_net),
            .ce(N__6567),
            .sr(N__6490));
    defparam o_X_1__nesr_3_LC_7_23_5.C_ON=1'b0;
    defparam o_X_1__nesr_3_LC_7_23_5.SEQ_MODE=4'b1000;
    defparam o_X_1__nesr_3_LC_7_23_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_1__nesr_3_LC_7_23_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3692),
            .lcout(o_X_c_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_1__nesr_3C_net),
            .ce(N__6568),
            .sr(N__6491));
    defparam o_X_1__nesr_5_LC_7_25_7.C_ON=1'b0;
    defparam o_X_1__nesr_5_LC_7_25_7.SEQ_MODE=4'b1000;
    defparam o_X_1__nesr_5_LC_7_25_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_1__nesr_5_LC_7_25_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4298),
            .lcout(o_X_c_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_1__nesr_5C_net),
            .ce(N__6569),
            .sr(N__6498));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_1_0_c_RNO_LC_9_18_0 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_1_0_c_RNO_LC_9_18_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_1_0_c_RNO_LC_9_18_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_1_0_c_RNO_LC_9_18_0  (
            .in0(N__5929),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_4_0_c_RNO_LC_9_18_1 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_4_0_c_RNO_LC_9_18_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_4_0_c_RNO_LC_9_18_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_4_0_c_RNO_LC_9_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5933),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_7_0_c_RNO_LC_9_18_2 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_7_0_c_RNO_LC_9_18_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_7_0_c_RNO_LC_9_18_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_7_0_c_RNO_LC_9_18_2  (
            .in0(N__5935),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_5_ma_LC_9_18_3 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_5_ma_LC_9_18_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_5_ma_LC_9_18_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_5_ma_LC_9_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5934),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_5_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_2_0_c_RNO_LC_9_18_4 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_2_0_c_RNO_LC_9_18_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_2_0_c_RNO_LC_9_18_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_2_0_c_RNO_LC_9_18_4  (
            .in0(N__5931),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_5_ma_LC_9_18_5 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_5_ma_LC_9_18_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_5_ma_LC_9_18_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_5_ma_LC_9_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5930),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_5_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_3_0_c_RNO_LC_9_18_6 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_3_0_c_RNO_LC_9_18_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_3_0_c_RNO_LC_9_18_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_3_0_c_RNO_LC_9_18_6  (
            .in0(N__5932),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_0_0_c_RNO_LC_9_18_7 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_0_0_c_RNO_LC_9_18_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_0_0_c_RNO_LC_9_18_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_0_0_c_RNO_LC_9_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5928),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_0_0_c_LC_9_19_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_0_0_c_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_0_0_c_LC_9_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_0_0_c_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3575),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_619 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_LUT4_0_LC_9_19_1 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_LUT4_0_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_LUT4_0_LC_9_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_LUT4_0_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3566),
            .in3(N__3557),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_619_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_619 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_620 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_620_THRU_LUT4_0_LC_9_19_2 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_620_THRU_LUT4_0_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_620_THRU_LUT4_0_LC_9_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_620_THRU_LUT4_0_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3554),
            .in3(N__3545),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_620_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_620 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_621 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_621_THRU_LUT4_0_LC_9_19_3 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_621_THRU_LUT4_0_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_621_THRU_LUT4_0_LC_9_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_621_THRU_LUT4_0_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3542),
            .in3(N__3533),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_621_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_621 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_622 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_622_THRU_LUT4_0_LC_9_19_4 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_622_THRU_LUT4_0_LC_9_19_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_622_THRU_LUT4_0_LC_9_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_622_THRU_LUT4_0_LC_9_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3632),
            .in3(N__3623),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_622_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_622 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_4_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_4_0_c_RNIHHTP_LC_9_19_5 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_4_0_c_RNIHHTP_LC_9_19_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_4_0_c_RNIHHTP_LC_9_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_4_0_c_RNIHHTP_LC_9_19_5  (
            .in0(_gnd_net_),
            .in1(N__6044),
            .in2(N__3620),
            .in3(N__3611),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_623 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_4_4 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_5_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_5_0_c_RNITTRA_LC_9_19_6 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_5_0_c_RNITTRA_LC_9_19_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_5_0_c_RNITTRA_LC_9_19_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_5_0_c_RNITTRA_LC_9_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5969),
            .in3(N__3608),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_624 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_5_4 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_625 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_625_THRU_LUT4_0_LC_9_19_7 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_625_THRU_LUT4_0_LC_9_19_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_625_THRU_LUT4_0_LC_9_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_625_THRU_LUT4_0_LC_9_19_7  (
            .in0(_gnd_net_),
            .in1(N__3605),
            .in2(_gnd_net_),
            .in3(N__3599),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_625_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_625 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_626 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_626_THRU_LUT4_0_LC_9_20_0 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_626_THRU_LUT4_0_LC_9_20_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_626_THRU_LUT4_0_LC_9_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_626_THRU_LUT4_0_LC_9_20_0  (
            .in0(_gnd_net_),
            .in1(N__3587),
            .in2(_gnd_net_),
            .in3(N__3596),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_626_THRU_CO ),
            .ltout(),
            .carryin(bfn_9_20_0_),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_627 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_627_THRU_LUT4_0_LC_9_20_1 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_627_THRU_LUT4_0_LC_9_20_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_627_THRU_LUT4_0_LC_9_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_627_THRU_LUT4_0_LC_9_20_1  (
            .in0(_gnd_net_),
            .in1(N__3581),
            .in2(_gnd_net_),
            .in3(N__3593),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_627_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_627 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_628 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_7_0_c_RNIVTM7_LC_9_20_2 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_7_0_c_RNIVTM7_LC_9_20_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_7_0_c_RNIVTM7_LC_9_20_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_7_0_c_RNIVTM7_LC_9_20_2  (
            .in0(_gnd_net_),
            .in1(N__4538),
            .in2(_gnd_net_),
            .in3(N__3590),
            .lcout(\DFT.multiplier.regsA_un3_result_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_8_0_c_RNO_LC_9_20_3 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_8_0_c_RNO_LC_9_20_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_8_0_c_RNO_LC_9_20_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_8_0_c_RNO_LC_9_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5952),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_9_0_c_RNO_LC_9_20_4 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_9_0_c_RNO_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_9_0_c_RNO_LC_9_20_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_9_0_c_RNO_LC_9_20_4  (
            .in0(N__5953),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.o_X_1__nesr_8_LC_9_22_0 .C_ON=1'b0;
    defparam \DFT.o_X_1__nesr_8_LC_9_22_0 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_1__nesr_8_LC_9_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_1__nesr_8_LC_9_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4633),
            .lcout(X_1__8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_1__nesr_8C_net ),
            .ce(N__4750),
            .sr(N__6495));
    defparam \DFT.o_X_1__nesr_7_LC_9_23_4 .C_ON=1'b0;
    defparam \DFT.o_X_1__nesr_7_LC_9_23_4 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_1__nesr_7_LC_9_23_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \DFT.o_X_1__nesr_7_LC_9_23_4  (
            .in0(_gnd_net_),
            .in1(N__4658),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(X_1__7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_1__nesr_7C_net ),
            .ce(N__4758),
            .sr(N__6499));
    defparam \DFT.o_X_1__nesr_9_LC_9_23_5 .C_ON=1'b0;
    defparam \DFT.o_X_1__nesr_9_LC_9_23_5 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_1__nesr_9_LC_9_23_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_1__nesr_9_LC_9_23_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4646),
            .lcout(X_1__9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_1__nesr_7C_net ),
            .ce(N__4758),
            .sr(N__6499));
    defparam o_X_1__nesr_1_LC_9_24_0.C_ON=1'b0;
    defparam o_X_1__nesr_1_LC_9_24_0.SEQ_MODE=4'b1000;
    defparam o_X_1__nesr_1_LC_9_24_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_1__nesr_1_LC_9_24_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3683),
            .lcout(o_X_c_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_1__nesr_1C_net),
            .ce(N__6571),
            .sr(N__6502));
    defparam o_X_1__nesr_7_LC_9_24_3.C_ON=1'b0;
    defparam o_X_1__nesr_7_LC_9_24_3.SEQ_MODE=4'b1000;
    defparam o_X_1__nesr_7_LC_9_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_1__nesr_7_LC_9_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4286),
            .lcout(o_X_c_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_1__nesr_1C_net),
            .ce(N__6571),
            .sr(N__6502));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_0_0_c_LC_10_17_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_0_0_c_LC_10_17_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_0_0_c_LC_10_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_0_0_c_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4472),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_17_0_),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_583 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_583_THRU_LUT4_0_LC_10_17_1 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_583_THRU_LUT4_0_LC_10_17_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_583_THRU_LUT4_0_LC_10_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_583_THRU_LUT4_0_LC_10_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3824),
            .in3(N__3641),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_583_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_583 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_584 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_584_THRU_LUT4_0_LC_10_17_2 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_584_THRU_LUT4_0_LC_10_17_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_584_THRU_LUT4_0_LC_10_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_584_THRU_LUT4_0_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3815),
            .in3(N__3638),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_584_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_584 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_585 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_585_THRU_LUT4_0_LC_10_17_3 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_585_THRU_LUT4_0_LC_10_17_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_585_THRU_LUT4_0_LC_10_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_585_THRU_LUT4_0_LC_10_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3833),
            .in3(N__3635),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_585_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_585 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_586 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_586_THRU_LUT4_0_LC_10_17_4 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_586_THRU_LUT4_0_LC_10_17_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_586_THRU_LUT4_0_LC_10_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_586_THRU_LUT4_0_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4856),
            .in3(N__3737),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_586_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_586 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_4_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_4_0_c_RNIGMTH_LC_10_17_5 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_4_0_c_RNIGMTH_LC_10_17_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_4_0_c_RNIGMTH_LC_10_17_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_4_0_c_RNIGMTH_LC_10_17_5  (
            .in0(_gnd_net_),
            .in1(N__5402),
            .in2(N__3734),
            .in3(N__3725),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_587 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_4_5 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_5_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_5_0_c_RNIS2SI_LC_10_17_6 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_5_0_c_RNIS2SI_LC_10_17_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_5_0_c_RNIS2SI_LC_10_17_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_5_0_c_RNIS2SI_LC_10_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5393),
            .in3(N__3722),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_588 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_5_5 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_589 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_589_THRU_LUT4_0_LC_10_17_7 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_589_THRU_LUT4_0_LC_10_17_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_589_THRU_LUT4_0_LC_10_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_589_THRU_LUT4_0_LC_10_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5414),
            .in3(N__3719),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_589_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_589 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_590 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_590_THRU_LUT4_0_LC_10_18_0 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_590_THRU_LUT4_0_LC_10_18_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_590_THRU_LUT4_0_LC_10_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_590_THRU_LUT4_0_LC_10_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5702),
            .in3(N__3716),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_590_THRU_CO ),
            .ltout(),
            .carryin(bfn_10_18_0_),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_591 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_591_THRU_LUT4_0_LC_10_18_1 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_591_THRU_LUT4_0_LC_10_18_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_591_THRU_LUT4_0_LC_10_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_591_THRU_LUT4_0_LC_10_18_1  (
            .in0(_gnd_net_),
            .in1(N__5510),
            .in2(_gnd_net_),
            .in3(N__3713),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_591_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_591 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_592 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_592_THRU_LUT4_0_LC_10_18_2 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_592_THRU_LUT4_0_LC_10_18_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_592_THRU_LUT4_0_LC_10_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_592_THRU_LUT4_0_LC_10_18_2  (
            .in0(_gnd_net_),
            .in1(N__5000),
            .in2(_gnd_net_),
            .in3(N__3710),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_592_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_592 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_593 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_593_THRU_LUT4_0_LC_10_18_3 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_593_THRU_LUT4_0_LC_10_18_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_593_THRU_LUT4_0_LC_10_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_593_THRU_LUT4_0_LC_10_18_3  (
            .in0(_gnd_net_),
            .in1(N__4670),
            .in2(_gnd_net_),
            .in3(N__3707),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_593_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_593 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_594 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_594_THRU_LUT4_0_LC_10_18_4 .C_ON=1'b0;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_594_THRU_LUT4_0_LC_10_18_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_594_THRU_LUT4_0_LC_10_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_594_THRU_LUT4_0_LC_10_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3704),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_594_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_3_0_c_RNO_LC_10_18_5 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_3_0_c_RNO_LC_10_18_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_3_0_c_RNO_LC_10_18_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_3_0_c_RNO_LC_10_18_5  (
            .in0(N__5927),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_1_0_c_RNO_LC_10_18_6 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_1_0_c_RNO_LC_10_18_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_1_0_c_RNO_LC_10_18_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_1_0_c_RNO_LC_10_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5925),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_2_0_c_RNO_LC_10_18_7 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_2_0_c_RNO_LC_10_18_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_2_0_c_RNO_LC_10_18_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_2_0_c_RNO_LC_10_18_7  (
            .in0(N__5926),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_2_c_LC_10_19_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_2_c_LC_10_19_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_2_c_LC_10_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_2_c_LC_10_19_0  (
            .in0(_gnd_net_),
            .in1(N__4244),
            .in2(N__3806),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_10_19_0_),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_2_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_3_c_LC_10_19_1 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_3_c_LC_10_19_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_3_c_LC_10_19_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_3_c_LC_10_19_1  (
            .in0(_gnd_net_),
            .in1(N__4403),
            .in2(N__3794),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_2_4 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_3_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIS12B1_LC_10_19_2 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIS12B1_LC_10_19_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIS12B1_LC_10_19_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIS12B1_LC_10_19_2  (
            .in0(_gnd_net_),
            .in1(N__4388),
            .in2(N__3782),
            .in3(N__3770),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_823 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_3_3 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_4_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNIK3NM_LC_10_19_3 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNIK3NM_LC_10_19_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNIK3NM_LC_10_19_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNIK3NM_LC_10_19_3  (
            .in0(_gnd_net_),
            .in1(N__4376),
            .in2(N__3767),
            .in3(N__3755),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_824 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_4_2 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_5_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIND4V_LC_10_19_4 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIND4V_LC_10_19_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIND4V_LC_10_19_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIND4V_LC_10_19_4  (
            .in0(_gnd_net_),
            .in1(N__4361),
            .in2(N__3752),
            .in3(N__3740),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_825 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_5_3 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_6_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNI50A41_LC_10_19_5 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNI50A41_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNI50A41_LC_10_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNI50A41_LC_10_19_5  (
            .in0(_gnd_net_),
            .in1(N__4349),
            .in2(N__3956),
            .in3(N__3944),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_826 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_6_1 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_7_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_7_c_RNINH451_LC_10_19_6 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_7_c_RNINH451_LC_10_19_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_7_c_RNINH451_LC_10_19_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_7_c_RNINH451_LC_10_19_6  (
            .in0(_gnd_net_),
            .in1(N__3941),
            .in2(N__4340),
            .in3(N__3932),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_827 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_7_1 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_8_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_8_c_RNIQRHD_LC_10_19_7 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_8_c_RNIQRHD_LC_10_19_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_8_c_RNIQRHD_LC_10_19_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_8_c_RNIQRHD_LC_10_19_7  (
            .in0(_gnd_net_),
            .in1(N__4328),
            .in2(N__3929),
            .in3(N__3920),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_828 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_8_1 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_9_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_9_c_RNI4O6E_LC_10_20_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_9_c_RNI4O6E_LC_10_20_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_9_c_RNI4O6E_LC_10_20_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_9_c_RNI4O6E_LC_10_20_0  (
            .in0(_gnd_net_),
            .in1(N__4313),
            .in2(N__3917),
            .in3(N__3905),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_829 ),
            .ltout(),
            .carryin(bfn_10_20_0_),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_10_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_10_c_RNIE7KN_LC_10_20_1 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_10_c_RNIE7KN_LC_10_20_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_10_c_RNIE7KN_LC_10_20_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_10_c_RNIE7KN_LC_10_20_1  (
            .in0(_gnd_net_),
            .in1(N__3902),
            .in2(N__4517),
            .in3(N__3893),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_830 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_10_0 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_11_c_RNIO44O_LC_10_20_2 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_11_c_RNIO44O_LC_10_20_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_11_c_RNIO44O_LC_10_20_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_11_c_RNIO44O_LC_10_20_2  (
            .in0(_gnd_net_),
            .in1(N__4502),
            .in2(N__3890),
            .in3(N__3878),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_831 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_11 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_12_c_RNIQFFJ1_LC_10_20_3 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_12_c_RNIQFFJ1_LC_10_20_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_12_c_RNIQFFJ1_LC_10_20_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_1_regsA_un3_result_cry_12_c_RNIQFFJ1_LC_10_20_3  (
            .in0(N__4481),
            .in1(N__3998),
            .in2(N__3875),
            .in3(N__3866),
            .lcout(\DFT.multiplier.regsA_un3_result_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_RNI8J5C1_LC_10_21_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_RNI8J5C1_LC_10_21_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_RNI8J5C1_LC_10_21_0 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_RNI8J5C1_LC_10_21_0  (
            .in0(N__4222),
            .in1(N__4462),
            .in2(N__3863),
            .in3(N__4463),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNI8J5C1 ),
            .ltout(),
            .carryin(bfn_10_21_0_),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_2_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_2_c_RNID4E01_LC_10_21_1 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_2_c_RNID4E01_LC_10_21_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_2_c_RNID4E01_LC_10_21_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_2_c_RNID4E01_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__4445),
            .in2(N__3848),
            .in3(N__3836),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_860 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_2_3 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_3_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_3_c_RNIMULJ1_LC_10_21_2 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_3_c_RNIMULJ1_LC_10_21_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_3_c_RNIMULJ1_LC_10_21_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_3_c_RNIMULJ1_LC_10_21_2  (
            .in0(_gnd_net_),
            .in1(N__4061),
            .in2(N__4433),
            .in3(N__4052),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_861 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_3_2 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_4_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_4_c_RNI4HRO_LC_10_21_3 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_4_c_RNI4HRO_LC_10_21_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_4_c_RNI4HRO_LC_10_21_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_4_c_RNI4HRO_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(N__4049),
            .in2(N__4418),
            .in3(N__4040),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_862 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_4_1 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_5_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_5_c_RNISIG41_LC_10_21_4 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_5_c_RNISIG41_LC_10_21_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_5_c_RNISIG41_LC_10_21_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_5_c_RNISIG41_LC_10_21_4  (
            .in0(_gnd_net_),
            .in1(N__4580),
            .in2(N__4037),
            .in3(N__4025),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_863 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_5_2 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_6_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_6_c_RNIA5M91_LC_10_21_5 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_6_c_RNIA5M91_LC_10_21_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_6_c_RNIA5M91_LC_10_21_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_6_c_RNIA5M91_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__4022),
            .in2(N__4568),
            .in3(N__4016),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_864 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_6_0 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_7_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_7_c_RNISMGA1_LC_10_21_6 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_7_c_RNISMGA1_LC_10_21_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_7_c_RNISMGA1_LC_10_21_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_2_regsA_un3_result_cry_7_c_RNISMGA1_LC_10_21_6  (
            .in0(_gnd_net_),
            .in1(N__4553),
            .in2(N__4013),
            .in3(N__4004),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_865 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_7_0 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.regsA_un3_result_cry_8_THRU_LUT4_0_LC_10_21_7 .C_ON=1'b0;
    defparam \DFT.multiplier.regsA_un3_result_cry_8_THRU_LUT4_0_LC_10_21_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.regsA_un3_result_cry_8_THRU_LUT4_0_LC_10_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.regsA_un3_result_cry_8_THRU_LUT4_0_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4001),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_8_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.o_X_1__nesr_6_LC_10_22_0 .C_ON=1'b1;
    defparam \DFT.o_X_1__nesr_6_LC_10_22_0 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_1__nesr_6_LC_10_22_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \DFT.o_X_1__nesr_6_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__5686),
            .in2(N__5662),
            .in3(_gnd_net_),
            .lcout(X_1__6),
            .ltout(),
            .carryin(bfn_10_22_0_),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_2_1 ),
            .clk(\INVDFT.o_X_1__nesr_6C_net ),
            .ce(N__4751),
            .sr(N__6496));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_2_c_RNIMU8V_LC_10_22_1 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_2_c_RNIMU8V_LC_10_22_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_2_c_RNIMU8V_LC_10_22_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_2_c_RNIMU8V_LC_10_22_1  (
            .in0(_gnd_net_),
            .in1(N__3983),
            .in2(N__3971),
            .in3(N__3959),
            .lcout(\DFT.x_7 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_2_1 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_3_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIQ8CH2_LC_10_22_2 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIQ8CH2_LC_10_22_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIQ8CH2_LC_10_22_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIQ8CH2_LC_10_22_2  (
            .in0(_gnd_net_),
            .in1(N__4229),
            .in2(N__4223),
            .in3(N__4205),
            .lcout(\DFT.x_8 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_3_0 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_4_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNIEERA2_LC_10_22_3 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNIEERA2_LC_10_22_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNIEERA2_LC_10_22_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNIEERA2_LC_10_22_3  (
            .in0(_gnd_net_),
            .in1(N__4202),
            .in2(N__4193),
            .in3(N__4184),
            .lcout(\DFT.x_9 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_4_8 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_5_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIASUU2_LC_10_22_4 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIASUU2_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIASUU2_LC_10_22_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIASUU2_LC_10_22_4  (
            .in0(_gnd_net_),
            .in1(N__4181),
            .in2(N__4172),
            .in3(N__4163),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_963 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_5_1 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNISQIC1_LC_10_22_5 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNISQIC1_LC_10_22_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNISQIC1_LC_10_22_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNISQIC1_LC_10_22_5  (
            .in0(_gnd_net_),
            .in1(N__4160),
            .in2(N__4151),
            .in3(N__4142),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_964 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_6 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_7_c_RNIVQTO1_LC_10_22_6 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_7_c_RNIVQTO1_LC_10_22_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_7_c_RNIVQTO1_LC_10_22_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_7_c_RNIVQTO1_LC_10_22_6  (
            .in0(_gnd_net_),
            .in1(N__4139),
            .in2(N__4130),
            .in3(N__4121),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_965 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_7 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_8_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_8_c_RNIOUH72_LC_10_22_7 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_8_c_RNIOUH72_LC_10_22_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_8_c_RNIOUH72_LC_10_22_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_8_c_RNIOUH72_LC_10_22_7  (
            .in0(_gnd_net_),
            .in1(N__4118),
            .in2(N__4109),
            .in3(N__4100),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_966 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_8_0 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_9_c_RNILFT82_LC_10_23_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_9_c_RNILFT82_LC_10_23_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_9_c_RNILFT82_LC_10_23_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_9_c_RNILFT82_LC_10_23_0  (
            .in0(_gnd_net_),
            .in1(N__4097),
            .in2(N__4088),
            .in3(N__4076),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_967 ),
            .ltout(),
            .carryin(bfn_10_23_0_),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_10_c_RNITHMQ2_LC_10_23_1 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_10_c_RNITHMQ2_LC_10_23_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_10_c_RNITHMQ2_LC_10_23_1 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_3_m1_forloop_1_1_regsA_un3_result_cry_10_c_RNITHMQ2_LC_10_23_1  (
            .in0(N__5378),
            .in1(N__4073),
            .in2(N__4619),
            .in3(N__4064),
            .lcout(\DFT.multiplier.regsA_un3_result_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.o_X_1__nesr_12_LC_10_24_3 .C_ON=1'b0;
    defparam \DFT.o_X_1__nesr_12_LC_10_24_3 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_1__nesr_12_LC_10_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_1__nesr_12_LC_10_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4694),
            .lcout(X_1__12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_1__nesr_12C_net ),
            .ce(N__4763),
            .sr(N__6503));
    defparam \DFT.o_X_1__nesr_11_LC_10_24_6 .C_ON=1'b0;
    defparam \DFT.o_X_1__nesr_11_LC_10_24_6 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_1__nesr_11_LC_10_24_6 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \DFT.o_X_1__nesr_11_LC_10_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5312),
            .in3(_gnd_net_),
            .lcout(X_1__11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_1__nesr_12C_net ),
            .ce(N__4763),
            .sr(N__6503));
    defparam \DFT.o_X_1__nesr_13_LC_10_24_7 .C_ON=1'b0;
    defparam \DFT.o_X_1__nesr_13_LC_10_24_7 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_1__nesr_13_LC_10_24_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_1__nesr_13_LC_10_24_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4706),
            .lcout(X_1__13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_1__nesr_12C_net ),
            .ce(N__4763),
            .sr(N__6503));
    defparam o_X_1__nesr_6_LC_10_25_5.C_ON=1'b0;
    defparam o_X_1__nesr_6_LC_10_25_5.SEQ_MODE=4'b1000;
    defparam o_X_1__nesr_6_LC_10_25_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_1__nesr_6_LC_10_25_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4280),
            .lcout(o_X_c_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_1__nesr_6C_net),
            .ce(N__6573),
            .sr(N__6507));
    defparam o_X_1__nesr_4_LC_10_26_6.C_ON=1'b0;
    defparam o_X_1__nesr_4_LC_10_26_6.SEQ_MODE=4'b1000;
    defparam o_X_1__nesr_4_LC_10_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_1__nesr_4_LC_10_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4604),
            .lcout(o_X_c_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_1__nesr_4C_net),
            .ce(N__6575),
            .sr(N__6511));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_0_0_c_LC_11_17_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_0_0_c_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_0_0_c_LC_11_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_0_0_c_LC_11_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4865),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_17_0_),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_1_0_c_LC_11_17_1 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_1_0_c_LC_11_17_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_1_0_c_LC_11_17_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_1_0_c_LC_11_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4874),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_0 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_2_0_c_LC_11_17_2 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_2_0_c_LC_11_17_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_2_0_c_LC_11_17_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_2_0_c_LC_11_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4892),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_1 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_549 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_549_THRU_LUT4_0_LC_11_17_3 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_549_THRU_LUT4_0_LC_11_17_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_549_THRU_LUT4_0_LC_11_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_549_THRU_LUT4_0_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4883),
            .in3(N__4232),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_549_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_549 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_550 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_550_THRU_LUT4_0_LC_11_17_4 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_550_THRU_LUT4_0_LC_11_17_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_550_THRU_LUT4_0_LC_11_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_550_THRU_LUT4_0_LC_11_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4829),
            .in3(N__4391),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_550_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_550 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_4_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_4_0_c_RNIQ3MM_LC_11_17_5 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_4_0_c_RNIQ3MM_LC_11_17_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_4_0_c_RNIQ3MM_LC_11_17_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_4_0_c_RNIQ3MM_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5018),
            .in3(N__4379),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_551 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_4_6 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_5_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_5_0_c_RNIGV3E_LC_11_17_6 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_5_0_c_RNIGV3E_LC_11_17_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_5_0_c_RNIGV3E_LC_11_17_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_5_0_c_RNIGV3E_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(N__4835),
            .in2(N__4844),
            .in3(N__4364),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_552 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_5_6 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_553 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_553_THRU_LUT4_0_LC_11_17_7 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_553_THRU_LUT4_0_LC_11_17_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_553_THRU_LUT4_0_LC_11_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_553_THRU_LUT4_0_LC_11_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5027),
            .in3(N__4352),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_553_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_553 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_554 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_554_THRU_LUT4_0_LC_11_18_0 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_554_THRU_LUT4_0_LC_11_18_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_554_THRU_LUT4_0_LC_11_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_554_THRU_LUT4_0_LC_11_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5036),
            .in3(N__4343),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_554_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_18_0_),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_555 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_555_THRU_LUT4_0_LC_11_18_1 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_555_THRU_LUT4_0_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_555_THRU_LUT4_0_LC_11_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_555_THRU_LUT4_0_LC_11_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5105),
            .in3(N__4331),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_555_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_555 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_556 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_556_THRU_LUT4_0_LC_11_18_2 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_556_THRU_LUT4_0_LC_11_18_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_556_THRU_LUT4_0_LC_11_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_556_THRU_LUT4_0_LC_11_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5009),
            .in3(N__4316),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_556_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_556 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_557 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_557_THRU_LUT4_0_LC_11_18_3 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_557_THRU_LUT4_0_LC_11_18_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_557_THRU_LUT4_0_LC_11_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_557_THRU_LUT4_0_LC_11_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5360),
            .in3(N__4301),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_557_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_557 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_558 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_558_THRU_LUT4_0_LC_11_18_4 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_558_THRU_LUT4_0_LC_11_18_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_558_THRU_LUT4_0_LC_11_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_558_THRU_LUT4_0_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(N__5522),
            .in2(_gnd_net_),
            .in3(N__4505),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_558_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_558 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_559 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_559_THRU_LUT4_0_LC_11_18_5 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_559_THRU_LUT4_0_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_559_THRU_LUT4_0_LC_11_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_559_THRU_LUT4_0_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__4529),
            .in2(_gnd_net_),
            .in3(N__4493),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_559_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_559 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_560 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_11_0_c_RNIHNIP_LC_11_18_6 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_11_0_c_RNIHNIP_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_11_0_c_RNIHNIP_LC_11_18_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_11_0_c_RNIHNIP_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__4490),
            .in2(_gnd_net_),
            .in3(N__4484),
            .lcout(\DFT.multiplier.regsA_un3_result_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_0_0_c_RNO_LC_11_18_7 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_0_0_c_RNO_LC_11_18_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_0_0_c_RNO_LC_11_18_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_0_0_c_RNO_LC_11_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5868),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_LC_11_19_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_LC_11_19_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_LC_11_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_LC_11_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5246),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_655 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_655_THRU_LUT4_0_LC_11_19_1 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_655_THRU_LUT4_0_LC_11_19_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_655_THRU_LUT4_0_LC_11_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_655_THRU_LUT4_0_LC_11_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5291),
            .in3(N__4448),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_655_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_655 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_656 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_656_THRU_LUT4_0_LC_11_19_2 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_656_THRU_LUT4_0_LC_11_19_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_656_THRU_LUT4_0_LC_11_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_656_THRU_LUT4_0_LC_11_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5282),
            .in3(N__4436),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_656_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_656 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_657 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_657_THRU_LUT4_0_LC_11_19_3 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_657_THRU_LUT4_0_LC_11_19_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_657_THRU_LUT4_0_LC_11_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_657_THRU_LUT4_0_LC_11_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5264),
            .in3(N__4421),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_657_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_657 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_658 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_658_THRU_LUT4_0_LC_11_19_4 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_658_THRU_LUT4_0_LC_11_19_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_658_THRU_LUT4_0_LC_11_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_658_THRU_LUT4_0_LC_11_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5255),
            .in3(N__4406),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_658_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_658 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_4_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_4_0_c_RNIICTH_LC_11_19_5 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_4_0_c_RNIICTH_LC_11_19_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_4_0_c_RNIICTH_LC_11_19_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_4_0_c_RNIICTH_LC_11_19_5  (
            .in0(_gnd_net_),
            .in1(N__4991),
            .in2(N__5273),
            .in3(N__4571),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_659 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_4_7 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_5_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_5_0_c_RNIUORI_LC_11_19_6 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_5_0_c_RNIUORI_LC_11_19_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_5_0_c_RNIUORI_LC_11_19_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_5_0_c_RNIUORI_LC_11_19_6  (
            .in0(_gnd_net_),
            .in1(N__5297),
            .in2(_gnd_net_),
            .in3(N__4556),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_660 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_5_7 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_661 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_661_THRU_LUT4_0_LC_11_19_7 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_661_THRU_LUT4_0_LC_11_19_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_661_THRU_LUT4_0_LC_11_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_661_THRU_LUT4_0_LC_11_19_7  (
            .in0(_gnd_net_),
            .in1(N__5498),
            .in2(_gnd_net_),
            .in3(N__4544),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_661_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_661 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_662 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_662_THRU_LUT4_0_LC_11_20_0 .C_ON=1'b0;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_662_THRU_LUT4_0_LC_11_20_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_662_THRU_LUT4_0_LC_11_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_662_THRU_LUT4_0_LC_11_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4541),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_662_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_13_0_c_RNO_LC_11_20_1 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_13_0_c_RNO_LC_11_20_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_13_0_c_RNO_LC_11_20_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_13_0_c_RNO_LC_11_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5944),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_13_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.state_RNIR1CE_0_LC_11_20_3 .C_ON=1'b0;
    defparam \DFT.state_RNIR1CE_0_LC_11_20_3 .SEQ_MODE=4'b0000;
    defparam \DFT.state_RNIR1CE_0_LC_11_20_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.state_RNIR1CE_0_LC_11_20_3  (
            .in0(N__5166),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5207),
            .lcout(\DFT.state_2_0 ),
            .ltout(\DFT.state_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.state_RNITIC91_1_LC_11_20_4 .C_ON=1'b0;
    defparam \DFT.state_RNITIC91_1_LC_11_20_4 .SEQ_MODE=4'b0000;
    defparam \DFT.state_RNITIC91_1_LC_11_20_4 .LUT_INIT=16'b1010111010101010;
    LogicCell40 \DFT.state_RNITIC91_1_LC_11_20_4  (
            .in0(N__6530),
            .in1(N__5167),
            .in2(N__4520),
            .in3(N__5065),
            .lcout(\DFT.un1_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.state_0_LC_11_20_5 .C_ON=1'b0;
    defparam \DFT.state_0_LC_11_20_5 .SEQ_MODE=4'b1000;
    defparam \DFT.state_0_LC_11_20_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \DFT.state_0_LC_11_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5091),
            .lcout(\DFT.stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.state_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.state_1_LC_11_20_6 .C_ON=1'b0;
    defparam \DFT.state_1_LC_11_20_6 .SEQ_MODE=4'b1000;
    defparam \DFT.state_1_LC_11_20_6 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \DFT.state_1_LC_11_20_6  (
            .in0(N__5092),
            .in1(N__5165),
            .in2(_gnd_net_),
            .in3(N__5066),
            .lcout(\DFT.stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.state_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_11_0_c_RNO_LC_11_20_7 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_11_0_c_RNO_LC_11_20_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_11_0_c_RNO_LC_11_20_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_11_0_c_RNO_LC_11_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5943),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.o_X_0__nesr_7_LC_11_21_1 .C_ON=1'b0;
    defparam \DFT.o_X_0__nesr_7_LC_11_21_1 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_0__nesr_7_LC_11_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_0__nesr_7_LC_11_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4657),
            .lcout(X_0__7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_0__nesr_7C_net ),
            .ce(N__5632),
            .sr(N__6497));
    defparam \DFT.o_X_0__nesr_9_LC_11_21_3 .C_ON=1'b0;
    defparam \DFT.o_X_0__nesr_9_LC_11_21_3 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_0__nesr_9_LC_11_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_0__nesr_9_LC_11_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4645),
            .lcout(X_0__9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_0__nesr_7C_net ),
            .ce(N__5632),
            .sr(N__6497));
    defparam \DFT.o_X_0__nesr_8_LC_11_21_5 .C_ON=1'b0;
    defparam \DFT.o_X_0__nesr_8_LC_11_21_5 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_0__nesr_8_LC_11_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_0__nesr_8_LC_11_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4634),
            .lcout(X_0__8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_0__nesr_7C_net ),
            .ce(N__5632),
            .sr(N__6497));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_RNIRG904_LC_11_22_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_RNIRG904_LC_11_22_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_RNIRG904_LC_11_22_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_RNIRG904_LC_11_22_0  (
            .in0(_gnd_net_),
            .in1(N__5237),
            .in2(N__5456),
            .in3(N__4789),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNIRG904 ),
            .ltout(),
            .carryin(bfn_11_22_0_),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.regsA_un3_result_cry_2_THRU_LUT4_0_LC_11_22_1 .C_ON=1'b0;
    defparam \DFT.multiplier.regsA_un3_result_cry_2_THRU_LUT4_0_LC_11_22_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.regsA_un3_result_cry_2_THRU_LUT4_0_LC_11_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.regsA_un3_result_cry_2_THRU_LUT4_0_LC_11_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4622),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.o_X_1__nesr_10_LC_11_23_0 .C_ON=1'b1;
    defparam \DFT.o_X_1__nesr_10_LC_11_23_0 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_1__nesr_10_LC_11_23_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \DFT.o_X_1__nesr_10_LC_11_23_0  (
            .in0(_gnd_net_),
            .in1(N__6143),
            .in2(N__5341),
            .in3(_gnd_net_),
            .lcout(X_1__10),
            .ltout(),
            .carryin(bfn_11_23_0_),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_2_0 ),
            .clk(\INVDFT.o_X_1__nesr_10C_net ),
            .ce(N__4762),
            .sr(N__6504));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_2_c_RNI1KHL1_LC_11_23_1 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_2_c_RNI1KHL1_LC_11_23_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_2_c_RNI1KHL1_LC_11_23_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_2_c_RNI1KHL1_LC_11_23_1  (
            .in0(_gnd_net_),
            .in1(N__6104),
            .in2(N__4592),
            .in3(N__4583),
            .lcout(\DFT.x_11 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_2_0 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIGSDC2_LC_11_23_2 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIGSDC2_LC_11_23_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIGSDC2_LC_11_23_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_3_c_RNIGSDC2_LC_11_23_2  (
            .in0(_gnd_net_),
            .in1(N__5489),
            .in2(N__4820),
            .in3(N__4811),
            .lcout(\DFT.x_12 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_3 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_4_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNI7QS33_LC_11_23_3 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNI7QS33_LC_11_23_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNI7QS33_LC_11_23_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_4_c_RNI7QS33_LC_11_23_3  (
            .in0(_gnd_net_),
            .in1(N__5474),
            .in2(N__4808),
            .in3(N__4799),
            .lcout(\DFT.x_13 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_4_0 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_5_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIEKOF6_LC_11_23_4 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIEKOF6_LC_11_23_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIEKOF6_LC_11_23_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_5_c_RNIEKOF6_LC_11_23_4  (
            .in0(_gnd_net_),
            .in1(N__4796),
            .in2(N__4790),
            .in3(N__4775),
            .lcout(\DFT.x_14 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_5_0 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_6_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNIS7913_LC_11_23_5 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNIS7913_LC_11_23_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNIS7913_LC_11_23_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_4_m1_forloop_1_1_regsA_un3_result_cry_6_c_RNIS7913_LC_11_23_5  (
            .in0(_gnd_net_),
            .in1(N__4772),
            .in2(_gnd_net_),
            .in3(N__4766),
            .lcout(\DFT.x_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.o_X_1__nesr_15_LC_11_23_6 .C_ON=1'b0;
    defparam \DFT.o_X_1__nesr_15_LC_11_23_6 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_1__nesr_15_LC_11_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_1__nesr_15_LC_11_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4681),
            .lcout(X_1__15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_1__nesr_10C_net ),
            .ce(N__4762),
            .sr(N__6504));
    defparam \DFT.o_X_1__nesr_14_LC_11_23_7 .C_ON=1'b0;
    defparam \DFT.o_X_1__nesr_14_LC_11_23_7 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_1__nesr_14_LC_11_23_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_1__nesr_14_LC_11_23_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5323),
            .lcout(X_1__14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_1__nesr_10C_net ),
            .ce(N__4762),
            .sr(N__6504));
    defparam \DFT.o_X_0__nesr_13_LC_11_24_3 .C_ON=1'b0;
    defparam \DFT.o_X_0__nesr_13_LC_11_24_3 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_0__nesr_13_LC_11_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_0__nesr_13_LC_11_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4705),
            .lcout(X_0__13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_0__nesr_13C_net ),
            .ce(N__5639),
            .sr(N__6508));
    defparam \DFT.o_X_0__nesr_12_LC_11_24_4 .C_ON=1'b0;
    defparam \DFT.o_X_0__nesr_12_LC_11_24_4 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_0__nesr_12_LC_11_24_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_0__nesr_12_LC_11_24_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4693),
            .lcout(X_0__12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_0__nesr_13C_net ),
            .ce(N__5639),
            .sr(N__6508));
    defparam \DFT.o_X_0__nesr_15_LC_11_24_6 .C_ON=1'b0;
    defparam \DFT.o_X_0__nesr_15_LC_11_24_6 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_0__nesr_15_LC_11_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_0__nesr_15_LC_11_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4682),
            .lcout(X_0__15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_0__nesr_13C_net ),
            .ce(N__5639),
            .sr(N__6508));
    defparam o_X_0__nesr_9_LC_11_26_4.C_ON=1'b0;
    defparam o_X_0__nesr_9_LC_11_26_4.SEQ_MODE=4'b1000;
    defparam o_X_0__nesr_9_LC_11_26_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_0__nesr_9_LC_11_26_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4985),
            .lcout(o_X_c_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_0__nesr_9C_net),
            .ce(N__6576),
            .sr(N__6513));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_2_0_c_RNO_LC_12_17_0 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_2_0_c_RNO_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_2_0_c_RNO_LC_12_17_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_2_0_c_RNO_LC_12_17_0  (
            .in0(N__5835),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_3_0_c_RNO_LC_12_17_1 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_3_0_c_RNO_LC_12_17_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_3_0_c_RNO_LC_12_17_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_3_0_c_RNO_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5836),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_1_0_c_RNO_LC_12_17_2 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_1_0_c_RNO_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_1_0_c_RNO_LC_12_17_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_1_0_c_RNO_LC_12_17_2  (
            .in0(N__5834),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_0_0_c_RNO_LC_12_17_3 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_0_0_c_RNO_LC_12_17_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_0_0_c_RNO_LC_12_17_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_0_0_c_RNO_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5833),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_4_0_c_RNO_LC_12_17_4 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_4_0_c_RNO_LC_12_17_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_4_0_c_RNO_LC_12_17_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_4_0_c_RNO_LC_12_17_4  (
            .in0(N__5837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_6_b_l_ofx_LC_12_17_5 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_6_b_l_ofx_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_6_b_l_ofx_LC_12_17_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_6_b_l_ofx_LC_12_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6032),
            .in3(N__5839),
            .lcout(\DFT.multiplier.regsA_un3_result_6_b_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_6_ma_LC_12_17_6 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_6_ma_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_6_ma_LC_12_17_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_6_ma_LC_12_17_6  (
            .in0(N__5840),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_6_ma_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_4_0_c_RNO_LC_12_17_7 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_4_0_c_RNO_LC_12_17_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_4_0_c_RNO_LC_12_17_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_4_0_c_RNO_LC_12_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5838),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.b_6_LC_12_18_0 .C_ON=1'b0;
    defparam \DFT.b_6_LC_12_18_0 .SEQ_MODE=4'b1000;
    defparam \DFT.b_6_LC_12_18_0 .LUT_INIT=16'b1000101011101010;
    LogicCell40 \DFT.b_6_LC_12_18_0  (
            .in0(N__6014),
            .in1(N__5221),
            .in2(N__5171),
            .in3(N__5077),
            .lcout(\DFT.bZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.b_6C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_9_0_c_RNO_LC_12_18_1 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_9_0_c_RNO_LC_12_18_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_9_0_c_RNO_LC_12_18_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_9_0_c_RNO_LC_12_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5876),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.a_0_LC_12_18_2 .C_ON=1'b0;
    defparam \DFT.a_0_LC_12_18_2 .SEQ_MODE=4'b1000;
    defparam \DFT.a_0_LC_12_18_2 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \DFT.a_0_LC_12_18_2  (
            .in0(N__5879),
            .in1(N__5096),
            .in2(_gnd_net_),
            .in3(N__5076),
            .lcout(\DFT.aZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.b_6C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_8_0_c_RNO_LC_12_18_3 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_8_0_c_RNO_LC_12_18_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_8_0_c_RNO_LC_12_18_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_8_0_c_RNO_LC_12_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5875),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_7_0_c_RNO_LC_12_18_4 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_7_0_c_RNO_LC_12_18_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_7_0_c_RNO_LC_12_18_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_7_0_c_RNO_LC_12_18_4  (
            .in0(N__5874),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_5_ma_LC_12_18_5 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_5_ma_LC_12_18_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_5_ma_LC_12_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_5_ma_LC_12_18_5  (
            .in0(_gnd_net_),
            .in1(N__5873),
            .in2(_gnd_net_),
            .in3(N__6013),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_5_ma_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_10_0_c_RNO_LC_12_18_6 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_10_0_c_RNO_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_10_0_c_RNO_LC_12_18_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_10_0_c_RNO_LC_12_18_6  (
            .in0(N__5877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_10_0_c_RNO_LC_12_18_7 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_10_0_c_RNO_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_10_0_c_RNO_LC_12_18_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_10_0_c_RNO_LC_12_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5878),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_10_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_5_b_l_ofx_LC_12_19_0 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_5_b_l_ofx_LC_12_19_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_5_b_l_ofx_LC_12_19_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_5_b_l_ofx_LC_12_19_0  (
            .in0(N__5885),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6026),
            .lcout(\DFT.multiplier.regsA_un3_result_5_b_l_ofx_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_6_ma_LC_12_19_1 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_6_ma_LC_12_19_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_6_ma_LC_12_19_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_6_ma_LC_12_19_1  (
            .in0(N__6027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5887),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_6_ma_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_1_0_c_RNO_LC_12_19_2 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_1_0_c_RNO_LC_12_19_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_1_0_c_RNO_LC_12_19_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_1_0_c_RNO_LC_12_19_2  (
            .in0(N__5881),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_2_0_c_RNO_LC_12_19_3 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_2_0_c_RNO_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_2_0_c_RNO_LC_12_19_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_2_0_c_RNO_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5882),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_5_ma_LC_12_19_4 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_5_ma_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_5_ma_LC_12_19_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_5_ma_LC_12_19_4  (
            .in0(N__5886),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_5_ma_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_3_0_c_RNO_LC_12_19_5 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_3_0_c_RNO_LC_12_19_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_3_0_c_RNO_LC_12_19_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_3_0_c_RNO_LC_12_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5883),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_4_0_c_RNO_LC_12_19_6 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_4_0_c_RNO_LC_12_19_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_4_0_c_RNO_LC_12_19_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_4_0_c_RNO_LC_12_19_6  (
            .in0(N__5884),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_RNO_LC_12_19_7 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_RNO_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_RNO_LC_12_19_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_0_0_c_RNO_LC_12_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5880),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_LC_12_20_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_LC_12_20_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_LC_12_20_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_LC_12_20_0  (
            .in0(_gnd_net_),
            .in1(N__5366),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_763 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_763_THRU_LUT4_0_LC_12_20_1 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_763_THRU_LUT4_0_LC_12_20_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_763_THRU_LUT4_0_LC_12_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_763_THRU_LUT4_0_LC_12_20_1  (
            .in0(_gnd_net_),
            .in1(N__5348),
            .in2(_gnd_net_),
            .in3(N__5225),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_763_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_763 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_764 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_1_0_c_RNIV67N_LC_12_20_2 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_1_0_c_RNIV67N_LC_12_20_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_1_0_c_RNIV67N_LC_12_20_2 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_1_0_c_RNIV67N_LC_12_20_2  (
            .in0(N__5423),
            .in1(N__5951),
            .in2(N__5954),
            .in3(N__5381),
            .lcout(\DFT.multiplier.regsA_un3_result_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_RNO_LC_12_20_3 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_RNO_LC_12_20_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_RNO_LC_12_20_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_0_0_c_RNO_LC_12_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5946),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_11_0_c_RNO_LC_12_20_5 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_11_0_c_RNO_LC_12_20_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_11_0_c_RNO_LC_12_20_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_11_0_c_RNO_LC_12_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5945),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_11_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_1_0_c_RNO_LC_12_20_6 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_1_0_c_RNO_LC_12_20_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_1_0_c_RNO_LC_12_20_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_7_regsA_un3_result_cry_1_0_c_RNO_LC_12_20_6  (
            .in0(N__5947),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.o_X_0__nesr_10_LC_12_22_0 .C_ON=1'b0;
    defparam \DFT.o_X_0__nesr_10_LC_12_22_0 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_0__nesr_10_LC_12_22_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DFT.o_X_0__nesr_10_LC_12_22_0  (
            .in0(_gnd_net_),
            .in1(N__6142),
            .in2(_gnd_net_),
            .in3(N__5342),
            .lcout(X_0__10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_0__nesr_10C_net ),
            .ce(N__5634),
            .sr(N__6505));
    defparam \DFT.o_X_0__nesr_14_LC_12_23_1 .C_ON=1'b0;
    defparam \DFT.o_X_0__nesr_14_LC_12_23_1 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_0__nesr_14_LC_12_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_0__nesr_14_LC_12_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5324),
            .lcout(X_0__14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_0__nesr_14C_net ),
            .ce(N__5633),
            .sr(N__6509));
    defparam \DFT.o_X_0__nesr_11_LC_12_24_6 .C_ON=1'b0;
    defparam \DFT.o_X_0__nesr_11_LC_12_24_6 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_0__nesr_11_LC_12_24_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.o_X_0__nesr_11_LC_12_24_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5308),
            .lcout(X_0__11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_0__nesr_11C_net ),
            .ce(N__5638),
            .sr(N__6512));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_6_a_LC_13_16_0 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_6_a_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_6_a_LC_13_16_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_6_a_LC_13_16_0  (
            .in0(N__5942),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6035),
            .lcout(\DFT.multiplier.regsA_un3_result_6_a ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_3_0_c_RNO_LC_13_16_1 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_3_0_c_RNO_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_3_0_c_RNO_LC_13_16_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_3_0_c_RNO_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5941),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_RNILH0D_LC_13_17_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_RNILH0D_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_RNILH0D_LC_13_17_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_RNILH0D_LC_13_17_0  (
            .in0(_gnd_net_),
            .in1(N__5531),
            .in2(N__6077),
            .in3(N__6076),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_897 ),
            .ltout(),
            .carryin(bfn_13_17_0_),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_2_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_2_c_RNII9QL_LC_13_17_1 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_2_c_RNII9QL_LC_13_17_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_2_c_RNII9QL_LC_13_17_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_2_c_RNII9QL_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(N__6053),
            .in2(N__6206),
            .in3(N__5459),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_898 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_2_2 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_3_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_3_c_RNIR3291_LC_13_17_2 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_3_c_RNIR3291_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_3_c_RNIR3291_LC_13_17_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_3_c_RNIR3291_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(N__6389),
            .in2(N__6188),
            .in3(N__5438),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_899 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_3_1 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_4_c_RNI9M7E_LC_13_17_3 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_4_c_RNI9M7E_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_4_c_RNI9M7E_LC_13_17_3 .LUT_INIT=16'b0110100110010110;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_2_m1_forloop_1_3_regsA_un3_result_cry_4_c_RNI9M7E_LC_13_17_3  (
            .in0(N__6170),
            .in1(N__6377),
            .in2(N__5435),
            .in3(N__5426),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_900 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_RNO_LC_13_17_4 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_RNO_LC_13_17_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_RNO_LC_13_17_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_RNO_LC_13_17_4  (
            .in0(N__5870),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_7_0_c_RNO_LC_13_17_5 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_7_0_c_RNO_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_7_0_c_RNO_LC_13_17_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_7_0_c_RNO_LC_13_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5872),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_5_b_l_ofx_LC_13_17_6 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_5_b_l_ofx_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_5_b_l_ofx_LC_13_17_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_5_b_l_ofx_LC_13_17_6  (
            .in0(N__5869),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6018),
            .lcout(\DFT.multiplier.regsA_un3_result_5_b_l_ofx_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_6_ma_LC_13_17_7 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_6_ma_LC_13_17_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_6_ma_LC_13_17_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_6_ma_LC_13_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6033),
            .in3(N__5871),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_6_ma_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_1_0_c_RNO_LC_13_18_0 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_1_0_c_RNO_LC_13_18_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_1_0_c_RNO_LC_13_18_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_1_0_c_RNO_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5889),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_3_0_c_RNO_LC_13_18_1 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_3_0_c_RNO_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_3_0_c_RNO_LC_13_18_1 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_3_0_c_RNO_LC_13_18_1  (
            .in0(N__5893),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_3_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_5_b_l_ofx_LC_13_18_2 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_5_b_l_ofx_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_5_b_l_ofx_LC_13_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_5_b_l_ofx_LC_13_18_2  (
            .in0(_gnd_net_),
            .in1(N__6028),
            .in2(_gnd_net_),
            .in3(N__5895),
            .lcout(\DFT.multiplier.regsA_un3_result_5_b_l_ofx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_1_0_c_RNO_LC_13_18_3 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_1_0_c_RNO_LC_13_18_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_1_0_c_RNO_LC_13_18_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_1_0_c_RNO_LC_13_18_3  (
            .in0(N__5890),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_1_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_0_0_c_RNO_LC_13_18_4 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_0_0_c_RNO_LC_13_18_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_0_0_c_RNO_LC_13_18_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_0_0_c_RNO_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5888),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_0_0_c_RNO_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_2_0_c_RNO_LC_13_18_5 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_2_0_c_RNO_LC_13_18_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_2_0_c_RNO_LC_13_18_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_2_0_c_RNO_LC_13_18_5  (
            .in0(N__5892),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_4_0_c_RNO_LC_13_18_6 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_4_0_c_RNO_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_4_0_c_RNO_LC_13_18_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_4_0_c_RNO_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5894),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_4_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_2_0_c_RNO_LC_13_18_7 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_2_0_c_RNO_LC_13_18_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_2_0_c_RNO_LC_13_18_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_2_0_c_RNO_LC_13_18_7  (
            .in0(N__5891),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_2_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_12_0_c_RNO_LC_13_19_0 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_12_0_c_RNO_LC_13_19_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_12_0_c_RNO_LC_13_19_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_1_regsA_un3_result_cry_12_0_c_RNO_LC_13_19_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5902),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_12_0_c_RNO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_9_0_c_RNO_LC_13_19_2 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_9_0_c_RNO_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_9_0_c_RNO_LC_13_19_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_9_0_c_RNO_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5899),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_9_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_7_0_c_RNO_LC_13_19_3 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_7_0_c_RNO_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_7_0_c_RNO_LC_13_19_3 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_4_regsA_un3_result_cry_7_0_c_RNO_LC_13_19_3  (
            .in0(N__5900),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_7_0_c_RNO_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_5_b_l_ofx_LC_13_19_4 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_5_b_l_ofx_LC_13_19_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_5_b_l_ofx_LC_13_19_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_5_b_l_ofx_LC_13_19_4  (
            .in0(_gnd_net_),
            .in1(N__5896),
            .in2(_gnd_net_),
            .in3(N__6022),
            .lcout(\DFT.multiplier.regsA_un3_result_5_b_l_ofx_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_6_ma_LC_13_19_5 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_6_ma_LC_13_19_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_6_ma_LC_13_19_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_3_regsA_un3_result_cry_6_ma_LC_13_19_5  (
            .in0(N__5897),
            .in1(_gnd_net_),
            .in2(N__6034),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_6_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_5_ma_LC_13_19_6 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_5_ma_LC_13_19_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_5_ma_LC_13_19_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_5_ma_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5901),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_5_ma ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_8_0_c_RNO_LC_13_19_7 .C_ON=1'b0;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_8_0_c_RNO_LC_13_19_7 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_8_0_c_RNO_LC_13_19_7 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_2_regsA_un3_result_cry_8_0_c_RNO_LC_13_19_7  (
            .in0(N__5898),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_8_0_c_RNO_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.o_X_0__nesr_6_LC_13_20_6 .C_ON=1'b0;
    defparam \DFT.o_X_0__nesr_6_LC_13_20_6 .SEQ_MODE=4'b1000;
    defparam \DFT.o_X_0__nesr_6_LC_13_20_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DFT.o_X_0__nesr_6_LC_13_20_6  (
            .in0(_gnd_net_),
            .in1(N__5687),
            .in2(_gnd_net_),
            .in3(N__5663),
            .lcout(X_0__6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVDFT.o_X_0__nesr_6C_net ),
            .ce(N__5622),
            .sr(N__6500));
    defparam o_X_0__nesr_7_LC_13_26_6.C_ON=1'b0;
    defparam o_X_0__nesr_7_LC_13_26_6.SEQ_MODE=4'b1000;
    defparam o_X_0__nesr_7_LC_13_26_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_0__nesr_7_LC_13_26_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5582),
            .lcout(o_X_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_0__nesr_7C_net),
            .ce(N__6580),
            .sr(N__6517));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_LC_14_17_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_LC_14_17_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_LC_14_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_6_regsA_un3_result_cry_0_0_c_LC_14_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5549),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_17_0_),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_727 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_727_THRU_LUT4_0_LC_14_17_1 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_727_THRU_LUT4_0_LC_14_17_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_727_THRU_LUT4_0_LC_14_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_727_THRU_LUT4_0_LC_14_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5540),
            .in3(N__5525),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_727_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_727 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_728 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_728_THRU_LUT4_0_LC_14_17_2 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_728_THRU_LUT4_0_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_728_THRU_LUT4_0_LC_14_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_728_THRU_LUT4_0_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__6212),
            .in2(_gnd_net_),
            .in3(N__6197),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_728_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_728 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_729 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_729_THRU_LUT4_0_LC_14_17_3 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_729_THRU_LUT4_0_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_729_THRU_LUT4_0_LC_14_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_729_THRU_LUT4_0_LC_14_17_3  (
            .in0(_gnd_net_),
            .in1(N__6194),
            .in2(_gnd_net_),
            .in3(N__6176),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_729_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_729 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_730 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_730_THRU_LUT4_0_LC_14_17_4 .C_ON=1'b0;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_730_THRU_LUT4_0_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_730_THRU_LUT4_0_LC_14_17_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_730_THRU_LUT4_0_LC_14_17_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6173),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_730_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_0_0_c_LC_14_18_0 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_0_0_c_LC_14_18_0 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_0_0_c_LC_14_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_0_0_c_LC_14_18_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6161),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_14_18_0_),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_691 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_LUT4_0_LC_14_18_1 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_LUT4_0_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_LUT4_0_LC_14_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_LUT4_0_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6152),
            .in3(N__6116),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_691_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_691 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_692 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_692_THRU_LUT4_0_LC_14_18_2 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_692_THRU_LUT4_0_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_692_THRU_LUT4_0_LC_14_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_692_THRU_LUT4_0_LC_14_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6113),
            .in3(N__6089),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_692_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_692 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_693 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_LUT4_0_LC_14_18_3 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_LUT4_0_LC_14_18_3 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_LUT4_0_LC_14_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_LUT4_0_LC_14_18_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6086),
            .in3(N__6062),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_693_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_693 ),
            .carryout(\DFT.multiplier.mult1_AdderTree2i_bigtree_694 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_694_THRU_LUT4_0_LC_14_18_4 .C_ON=1'b1;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_694_THRU_LUT4_0_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.mult1_AdderTree2i_bigtree_694_THRU_LUT4_0_LC_14_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.mult1_AdderTree2i_bigtree_694_THRU_LUT4_0_LC_14_18_4  (
            .in0(_gnd_net_),
            .in1(N__6059),
            .in2(_gnd_net_),
            .in3(N__6047),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_694_THRU_CO ),
            .ltout(),
            .carryin(\DFT.multiplier.mult1_AdderTree2i_bigtree_694 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_4_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_4_0_c_RNIJ7TP_LC_14_18_5 .C_ON=1'b1;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_4_0_c_RNIJ7TP_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_4_0_c_RNIJ7TP_LC_14_18_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \DFT.multiplier.o_x_if_w3_mult1_AdderTree2i_if_keep_adderTree_forloop2_1_m1_forloop_1_5_regsA_un3_result_cry_4_0_c_RNIJ7TP_LC_14_18_5  (
            .in0(_gnd_net_),
            .in1(N__6404),
            .in2(N__6398),
            .in3(N__6383),
            .lcout(\DFT.multiplier.mult1_AdderTree2i_bigtree_695 ),
            .ltout(),
            .carryin(\DFT.multiplier.regsA_un3_result_cry_4_3 ),
            .carryout(\DFT.multiplier.regsA_un3_result_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DFT.multiplier.regsA_un3_result_cry_5_THRU_LUT4_0_LC_14_18_6 .C_ON=1'b0;
    defparam \DFT.multiplier.regsA_un3_result_cry_5_THRU_LUT4_0_LC_14_18_6 .SEQ_MODE=4'b0000;
    defparam \DFT.multiplier.regsA_un3_result_cry_5_THRU_LUT4_0_LC_14_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DFT.multiplier.regsA_un3_result_cry_5_THRU_LUT4_0_LC_14_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6380),
            .lcout(\DFT.multiplier.regsA_un3_result_cry_5_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam o_X_0__nesr_1_LC_14_19_2.C_ON=1'b0;
    defparam o_X_0__nesr_1_LC_14_19_2.SEQ_MODE=4'b1000;
    defparam o_X_0__nesr_1_LC_14_19_2.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_0__nesr_1_LC_14_19_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6371),
            .lcout(o_X_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_0__nesr_1C_net),
            .ce(N__6570),
            .sr(N__6501));
    defparam o_X_0__nesr_0_LC_14_19_4.C_ON=1'b0;
    defparam o_X_0__nesr_0_LC_14_19_4.SEQ_MODE=4'b1000;
    defparam o_X_0__nesr_0_LC_14_19_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_0__nesr_0_LC_14_19_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6338),
            .lcout(o_X_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_0__nesr_1C_net),
            .ce(N__6570),
            .sr(N__6501));
    defparam o_X_1__nesr_8_LC_14_20_4.C_ON=1'b0;
    defparam o_X_1__nesr_8_LC_14_20_4.SEQ_MODE=4'b1000;
    defparam o_X_1__nesr_8_LC_14_20_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_1__nesr_8_LC_14_20_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6311),
            .lcout(o_X_c_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_1__nesr_8C_net),
            .ce(N__6572),
            .sr(N__6506));
    defparam o_X_0__nesr_3_LC_14_21_0.C_ON=1'b0;
    defparam o_X_0__nesr_3_LC_14_21_0.SEQ_MODE=4'b1000;
    defparam o_X_0__nesr_3_LC_14_21_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_0__nesr_3_LC_14_21_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6278),
            .lcout(o_X_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_0__nesr_3C_net),
            .ce(N__6574),
            .sr(N__6510));
    defparam o_X_0__nesr_2_LC_14_21_7.C_ON=1'b0;
    defparam o_X_0__nesr_2_LC_14_21_7.SEQ_MODE=4'b1000;
    defparam o_X_0__nesr_2_LC_14_21_7.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_0__nesr_2_LC_14_21_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6257),
            .lcout(o_X_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_0__nesr_3C_net),
            .ce(N__6574),
            .sr(N__6510));
    defparam o_X_0__nesr_4_LC_14_23_0.C_ON=1'b0;
    defparam o_X_0__nesr_4_LC_14_23_0.SEQ_MODE=4'b1000;
    defparam o_X_0__nesr_4_LC_14_23_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_0__nesr_4_LC_14_23_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6236),
            .lcout(o_X_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_0__nesr_4C_net),
            .ce(N__6577),
            .sr(N__6514));
    defparam o_X_0__nesr_8_LC_14_24_1.C_ON=1'b0;
    defparam o_X_0__nesr_8_LC_14_24_1.SEQ_MODE=4'b1000;
    defparam o_X_0__nesr_8_LC_14_24_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_0__nesr_8_LC_14_24_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6743),
            .lcout(o_X_c_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_0__nesr_8C_net),
            .ce(N__6579),
            .sr(N__6516));
    defparam o_X_1__nesr_9_LC_15_22_1.C_ON=1'b0;
    defparam o_X_1__nesr_9_LC_15_22_1.SEQ_MODE=4'b1000;
    defparam o_X_1__nesr_9_LC_15_22_1.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_1__nesr_9_LC_15_22_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6710),
            .lcout(o_X_c_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_1__nesr_9C_net),
            .ce(N__6578),
            .sr(N__6515));
    defparam o_X_0__nesr_5_LC_15_24_3.C_ON=1'b0;
    defparam o_X_0__nesr_5_LC_15_24_3.SEQ_MODE=4'b1000;
    defparam o_X_0__nesr_5_LC_15_24_3.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_0__nesr_5_LC_15_24_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6629),
            .lcout(o_X_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_0__nesr_5C_net),
            .ce(N__6581),
            .sr(N__6518));
    defparam o_X_0__nesr_6_LC_15_24_4.C_ON=1'b0;
    defparam o_X_0__nesr_6_LC_15_24_4.SEQ_MODE=4'b1000;
    defparam o_X_0__nesr_6_LC_15_24_4.LUT_INIT=16'b1111111100000000;
    LogicCell40 o_X_0__nesr_6_LC_15_24_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__6605),
            .lcout(o_X_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(INVo_X_0__nesr_5C_net),
            .ce(N__6581),
            .sr(N__6518));
    defparam CONSTANT_ONE_LUT4_LC_16_32_7.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_16_32_7.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_16_32_7.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_16_32_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // top_test
